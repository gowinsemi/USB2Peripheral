`protect begin_protected
`protect version="2.1"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2021-10",key_method="rsa"
`protect key_block
hVPVosDH2VwkuRZeYcJ2Tulh3wE2nb87TDmJh1/hn51uAlwq726GdEZYo/OS0T4jPrP60x6AEwMB
dDV5DFNWLLjgenCHitZNzFZZVVHKVjodGIr4WjWbzEqOQowonezzrWyaI1SkDRgSdGUOHvq58jV7
DIVPcceWM08BAu5ulbhtuSP6O7HIJko6j0xAy0WE1eKt70kb5TEQbhVvNPlNowVj52NrdeCy+YzR
HchwolxVeuqYnIMa7q7AatJ9NH9diOLc0+pYV2+VOHwykRrOdhsMzpZOsO4nafJ0nTu6bwUWR7Uo
7NWSG376Wg/ljm2tQZO80mU/XdKvQvVIqYQB7w==

`protect encoding=(enctype="base64", line_length=76, bytes=19504)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
HqPM1xGGK9zfxq/EAwBPQL8L8QcE6VbVaVAnLP8Q7zywVcohPXqdIP4wTtxaFbWRjuf464MzCTEc
bBkusM3lAqOSyhibRoS5vUhNMjEU+GDiRRF8BOKPbBBLl1i6dcni0JSCRCDIza+rCEFpEVls7jDe
PIVZ/XAkIq/dHJZKoKaAyWmCh/nLCh4tFnYtJhJiYTbk4B4hNizEx+P9xYaUPOS4b5R8jlwDzZsy
6BMTVBq7YkXOfQt3BEftxBbmbnsVMLlTYnk8zXzDqdohs0SGPgxuxKEjMAR3ugOdVH2bNcu3Lzbh
z1Vbvt6H84CCc8EZ88OatoZyinT9TNADPyxeF48u1lDo2741kx9BeYwvvSZadRxnz5/YAPqCcYM1
wbmx4UBQ8D/5unGd/Uu6b1MJlIPbTV06UrC8ekpVwJpp5EAfewEVahMzc4OpSAqgbjHqPcuKwHkf
hntxls7lffW5SAaREIDhxgCcAAO1BVZOGzjr7oXHzSS8gdP63XaU45jY8ON3LZaKEt0hEk87QVqn
qPQizkOEiOqjTQ4HoWwU8guxQTgu2PJBH1s3yd7Ot9mRGlQcGtzvxR6zBQrfU0VRpzde7Us54HEa
xYn5snfvXTVAETOrKxL4gD/f2wpribiohVCbH2NSEDeGpls76oskeVkF9oCOrfEH9PIpupWaNHis
MluTJ4hLzjQOYgqHFRIXgvCLSjTGFYcZD62LPgR1uAMC0KdlRE+9Z9GxLRpIK/YItVcig9IljO0z
2FbMy3IVZK6b/oT/U0wnaAIBCwkEitbytGk03yxNQzNPKQwG5hCPkn7gsBdj2cj53qEjsQMzYzcH
sM1+uvhXElDfKFk4ofguYYutUtGGF831InqjS5EwEMXL5dEcbUTASfE6y1q3SNx9J5pwRKsx6wjt
fFViiI0fO0yqqzwF8xn4BibT51S+Fmyky/g12tqo1BXv070+dU95vOK7VdSVXfYl1OFcz2NXuNj3
r//RnH6xN3e/gtmqH/BAG5gPdTxVkNuDBTyQGNpylbWGBkbqTLcHINSrNN5FEw9OeNUeIp1lcGpN
KjP5UROZ+w0EVQjaVfcCF2Ov+qF+8CEyJi1aSridTHyaITf2VAnU+kCxzusfon1mKUcR8OkwmLsA
sU9rGqJ65XbtZMGAFFb35rGe2cKo/K5oarxwyZ/+E78BBTZ3ZzN1HsdcSG65Q4rsrMXCTZ4U2OaG
fKSoGhpX7PYsymuX4rYtN3FR3KodRVJ5y2X2OmYWytZ50y0PliUYUpSVDCfH56lyK+mT74HRmzmj
ep+040/1EzyXXgb83XItw8JikOZAGuexDerMlRqe5ju72l+cdqHV/iE2ie+oBwg3b4yyIZISJUS1
l28pn2LHbIM/6CrXX3njkfEBSND1+syz+YUlCu50pvBYkIQuduUGNA8ZnvThwiaceHXj6kXzE26f
AEoMdjrRFAFCuBGa70vBEwEMYh1R698qtqSP/rJU3cjVrmGfQN72ukThlwNKycwRf6tgrTihriYD
17o3ETD9600dZDGAUuK9rZqpf/P5SKXzHacY/K3u0ULnJVb4CMLxfp6j0/5efxoDJrstxTUkY+X0
T51t87VNJ64CeCQ6dh1IuWI1VTFjsOO3rvJU8fi6qBBpq+Q/wKnKwvL+CJ9TkuNrWqmSXk6FUFVm
oeZLvDtdAQJrsrRE6E62i1wi4NSPKDw2maFFSu4hYFRQ6dmSGdKly6yvhHpCjvgI/BRCZg9Un77s
ndL/932NPBK0Pa/KWFjMXoBDIC+1DX2nuELZtsJnbCk+fYY/KRPRVX4PyMNQXloH1V5GnPZtlCyq
G3L38+2Te2G78AGfmsaGBEQKN6+NGLnrdNP6ZezpwWI9fNwvDDMKjN7BDJ/5+G35q1d72aJ8QR2z
zYZ/nHnx55r6Mj2Xz+fNBvkpm1siDPTH0l3oR61Z6+gEzs/7acpkZndDd6ZnzrYFOyCC9jFUCvYE
I7NIeTzO0iMTWuyVDCg209ZKwDZ89MRjwWPXkxotzhfYZJHYO2kmCMuPPJGlgR4nFxxwP71kxyHH
VF8JvLZSNLSEw2YmPOoshLptiuLvx9dDPCrCU273g3Dokeyb4un76eMmWNm/B4XdYAXl5VsXa5du
cE9OJZ4K6BxM8pvsq8sGbsm5UYoxD1CWmburmHMWIlodHRBHftmEMrEaVfzOtnlv+Q1qmUbBlqSO
pXGNSydZzrHOkj7ATT15JYLn3rsG1VM/ubDoHKOEgtjxRylhnT9aoQQJcrxriVuZBybK51iRWW4o
MdrXGQk871W9aJiWUbyOiw1dCF6TVQn5lXBK6lp4KztZXzNn5yIUgfgemp2Pk7RckzjclGuTtyGy
kc5FYEoj5XBNUk4As+NljfZkL1enqBoGA6FsBoV1frkWNlEHMFjfjWs67QOqJ9i63/Jj4GsGQb54
NHEyzXXn0vnUQ4b61IyopQTdu3k65h0Od5V47chiDxMlUhzlD6MUUYgf3HMWygUgXjg1pIOtIlE4
/cbm0XAnthaX9egokmtksmBYNz1JL3voxgPIviv2OE6R512Yidx5gXPlEwyJZunTK04ya233QXpi
T64FXWxlxgStnXufCEKItRRJ/g00RD9l+YnNa6Io//Vz4Jxh1Uqoq5qPBYthCvExWB6A/j1FSzox
w6AGJrMRqO+qxLATD6KhxA5a0OI5NHBEFabpuiCl7khXpya89Lg9E8PxrUzu0U0L4PV4Lx1jCKLS
63C+UgYbDbCmo0PXmoO+hgYsm/XDVCMSZI/YjJldRk8dPdZS5VT96K+27WYbP9+qgq7SjTDOOhAO
nfQKXGWCFWOqkMRezuRANUXHj9+7v+SlfdWANX6R3d8w1WDTo9pCk1Hy2lHGlArIg2j83KxVeXhp
JjGttU/+vZ5i80nstjwzON0wmJQhWvE2Fu2QfxcZRCVHHk/rGUYK9vzw54NxRYsRosPV2OsQISRn
A4dj3FjWOOrvlreSHi2fTAlzPyzQk6UFf6dPbZRTBY41qtjIjbJe+fW1nk9+p5dxf64F8r+5pGW3
dx4i42/jwLzPjR3CohNbsWHc72gvCRATEWecp6mxNDX+SmsZBO7omI+lqZM3MrLLhzPK+e+Tjwiu
AS4KD5R9Lwq4885jgECcb7aU+MFX9KD+BBCzffwrDpM/KJLJnS0eYgXmocNmPqUeWXPKIwq1RvLw
B7UWU/wYwEJ0rgw76uDucqoVAVYGTCzoezB6s8R58ZPUsWGxOIsgs2BR+udAztybpPkXoBRRcD30
AxcpAZ7O6bYP6J/WiMIKbl0i6taq7DyN7tudX18npdicfIDkBPtvoauahh4KjouSr0APwUkEk2tP
MuaXQRtMcgjPmeYA0doajf1QkK9xg5PBMKdz/uNa8sj4F9ZipTHO3WLI7ng49yuhlWJ/WQUvMIN5
QRplUfWE7tDH7eAOqA/Fr8T5Pq9BAtbRbfxh1VPt120OnYkqtFmyfNFv4Sj7wIrkPJCiUosuAZXW
/TwIve+Wuw/rqn3B0snTe9SwzYXK1R/3TwvSkS889vXeS9/HrFj7yVXxhqRU4f+IbzN4MnuESRSF
5oNnnoxpqeQloz9RHaNKXng0kQMs3msVwplfRuspzWfP4JD58pmUlcutkX1NvJui5iM5ETnwtfpb
DBIUHnetmHEx9bfPBpJSoeEqD+eMIN3fxLRT85iIBcTZgQ7PbQ6hHDK4IoardPW1FNrNgbKyNr9j
QZWmkXHufsaftGQq1+DwPpl3q3mMpwzC7rkrDLrQj3ZS2p9/JpoORYW0vf+tzTl/X9UeoZYiL2RN
kJDmdKZmchn6rR1d1ze5h0BignCNEDGYCF0NhEyAp/g7yBJCx7LHh5N70Kuan8vlsOLJM6UfmIfD
AhPa1cO1B6Q9qv+qrkvK2nQKFlTlIpKhx347cOwg3kD0VuMuQpn1KsbibFhAOkWHt6GK/rupUwa4
qZ0weZUqWUw9OoL222yLUiX4nTxb4Ejlp0ULh7ZWPgY5RgQaNR+tLUJTf+3AOd6342WJ5E4dvjbF
5zBrWJrMeFOdeiYB9qwOuDGCsTlWsP3a0QRJTePfuYwv/9v9b01TfvQ2cjnPgjQ/ewJRvon9gQHd
Ga48lNzAG9ieDqGx7GDiyuG6+hEVs+kfEUqfo1DPNmBzsZ2m7NpnzqWBIeWUBDZ70QXzGQX+dbzI
ao5q66m6RzJUoRmjbrmT3wLrFlRDgd+/hxDln+ic7jV1AJfpsHJOdOSg+vFuBCx+rqVE6Cbz2EXf
5riyefQqgTraqsxjDlkn/161VaL5ei3sD6JqvWp6wc1FDcjjl5j1jht8Rq11p6gGqnJbPyBmvbTN
anGE9mQ/wsM/S1TD3vly+mGubd+mJXlDdh6iIcHJ7jVrIrBdXme3bDgYLCdY2LqPQqvKQmE+Rv+P
IBeVJGDBeenN2GqOUOqwoPZdmxya07supBfmafH9QeY9lY7Vkd6x7g8ccm+piaXpHmc3YDz1mO0H
pyNvYayAfaOjdtuRT3WvXUvEfVL8scRVEsWOf22chni/MvCGtWjT1o7ypkhQqxmM6k8hnVsD4u70
+Zzq0n1EV+Xo7XxeeS51t3JFXO4E76/FwLIY65qL/sQlomcgRcpk/AXdDcJipmpRW8GefmD+R0UJ
PtD05tmH0UCdSEUtuSwIsFF7c9pSaMZQvHDZ43rTeNe9kECXAcfLZ6DVyYUN9u417N6w1Cbv7LCx
RrQeB78bMb+SItJdBX/ixpSMqBS35sAnfkIDadkF770GYAY9JtRJ9GcJsazN+T+ObFiSTezhcCKo
ZI2gE0444mtfeefEcfY4DA9cGLGRpA0HZaVVjf3+HfX+b0MfvkwMxBZtPXLkulHN/xifOrXbzXzs
wJqxKFozKeXYHXdY8X+WhNkJWZ6QPa0c2kGRXr7Y+PhdIsTl0/YI54+Ki87EKs/BJ6O4LkIdRO8Y
uXkSQ/bMVSMA7nxVvt7J/nwzd0qOpnJr8aUmC5aMIVazORgroCXnOZBP6EYTmiHzpF4oTEiV2xdE
StHqcbwh96VJsBojnTA7DSzSam7q4NOzHaG05apOY1icB/uCux//wiiWVHKPwpNalmekUhC1hi1C
IvoM8YfpSHm/J8kVQzN8LhK4yHZikXAZmoY6yjAS4lMEK0fR7Rrwx8QzlWHTbFdhHOckDWeRnmsi
9iMg7oahKXckIPz/dgnFUn3QJtqg9ZRpCEhshTvu2sY6w2IvRhjorLEmzpURTH+T815esTomIDkq
h2pMzwDQcKFHLEKv0MclILTEJs+lf7K4rNYeVWfTYYWjo+WTQ1zC0u9Krmkf06f2IDj88HvbtBiP
kjaZr0eo1zzTivklBCcpP4E2CTZH7XtZmSb9onci4cCoW3/bB1lxFtFDiXmCUifu4Y/7vZsjlOgD
udqzejAEmsrPLEm2fJnM7tVdkMCXSmG5Z11SN3BmtKt1aYIpJGANKLuwfKdSlqKFCwKZ0+Cr19Rx
WlfYc5QicoE7lUjeV+b0G6p7lIsYRrZ382cr02GHcNf2ecF1RemnMzWxtUB3C/vVQmT+Y+7GN9rT
mXijA0u01WsSYl9mKuGSB8Uav+KLAQYOe2g9jyjby50TNjI9/xkhW25pGRtgaoHVjiOEAeONyLoe
YzBmCmC+PIpf4bPC6Kj32cQIC3O7VbiKxXvTflp+xcFyFQEw7Ml4nQo92lt4OPX+5rrUjOCDu3Df
zjXf7YhTjn5BM/xM4BvVUwTb0B1OX6V+LPTOEjyDC3iX/aikn2QPkOs1Udra7UvBlOv5E4Gs/nq0
gsyfi/crvsBKkotgMibngjSJla0RN5B5oTpQU6+OLzyMRLnKnjPnGO/fv8n6YSeCzWLr/LFlOTim
8prfjNKIFrw/za/YSgk1rGu7ZqRyfoIFqNupueLR6LiL1GumIhVeOTF1seJZqfpC0B9E6OKCdmRW
JMtxo/eNfjgKQ6SuFM7XDo+YeHHNFKOEVdq1Txuoy2EjG6+yiYSw/+sY7aOG481nG02La5nv+z5g
Ysc32znR7ELyNWu2JSWlfxxqMiD7RGdHEIqOWDoXqWdOylYwDQ5cyDqPOnSyRTFWwszprNBT2hvk
wOt+ypmbFAazXIB68Gsu/zKFWk6d1fcNIW4pg4ASkndjUhLE2DxDqV+sK28RLqDAsiI7bW1xDeCP
VYDmqV0LzAS7o2LogBxm6P0AKfN1PuiQd9utaf7+UYWe6KwZxI5R7t59ffWjLYtEUuwBMng+xVJu
T0lQjOtNWXk1GGcxQhYxm2PzJcDCEiq+NehkNU9Aviz941IqfyYByvALX5jSXx/FmpWtJutjI0gy
G6h8z4Kg8S3op5N3b54wTGSuuLO44Qg60eP2ILe051fSJlBoGyLEAT3wzPDBv17OOrXao99O9Tqy
rJVeG3QEIjys8R3YrfHyxeDAi58AH83Ijmqt4Op3lC3RDI/aSITF9++ZIuPHVP16ZBfVEIAg536S
y3gm74xwxrFH2mxmbnb1fZUq7b1Mu/0pDjD0PPBPwhQhHnMxyZ7asHFlTQrIQRtJApucoo+qQAo+
Gm9Q3T5Z1dUAyslgV6+9C1SY0nuXofy9Lv63Ja302UVNDkU0yl0JWtSg6ZcmBwkUBATdTndw20eM
wjIlsB5GKVMdARPGj2mHEed3DiJdutd726+BL3TTFeDXK4GDj9tge+GDoXJ3++IwGmvesC0+HERs
2g5HIwZUoKEwQaALysBMhwFTzQqOAI1gXsLXb15QyjC3/O5cosa6OXmNFkGFJVFUQmipB1/YWdTn
da/U8an4zDuXAQg72tAr43k1fCeVtran/mCZCjG/LyGzyUX9mGaCCAcyqOJKkuV63BTtKMXuz15F
UcNX2LTg0orbAXCNxoyYsyCbj4FfaIc+X38lZjCBwGn4MsVgBBjTPxG+Bza8fqknwjOh7X3ND32N
MkEDBlpqt6EAZTCI09F8GnbELtcoYWZ5PG8e8sD5lbFew/DMlKari+pUg48U5atCybV+3c+OHwT0
lZkM1HlcAiivzzp2mg3F/Gfu/+JjSiwkOSg5Ii0gSI2C/18yotjp5Z/LAQ0m/SHEwOR3Le89j2Fg
L74skLZ2Z3gVieX4FePw6ylOF79PND8B5QnJHRL93OIwT2XWljguR0tIAZUO1Q/6d4LORCcJ/Qps
rrwLH2Eh9hbu+Aw0DjvaFZyAdlCMSEIvh8pNpw/2rvZC+N3Yuk6+C+3YdKf72eUQWoqmzbJjfmW7
n4Ne1LkpH9jsfDaV7BKYHhinfGTOYcpEttLSAcGw4gJtqrmcjrJmRTMzqlFkJuTnNspYgQTS2v4e
Rgptw36G86rcQr+jx1wGgzf77qCKhECshj2Ht3OArkcvl99SjXCet+rH7ZcTwhyp0VTaOcG/y48s
/cAEuFPjOjDpT+W9yE7QrdKLVpFflfQCd+WrKsPt0tYQid+HW1INnWKyfBVVdcHkGPHhz+hxmw9E
AOwGKhzm7n33046tPdQvVcxlXeFz7FuObPrffs3AClbAVRD+q1Xrg6gYoQ1alOjhFpJZ/rrDQDfb
+SkygX8N/fpARRCuznQAk8+npre7P8Kr1AA7PSoUu4dMKF11k3s99aznn/xcDbg3eHyOnnHxkDrI
vGA9NEr3/G2luXVXvXeWYznaFzTF71kFpr6886BHgqmYqf4nsa4Gbsi1riK6niwirgDP4YBbGDel
kxh1359KqLNiw5YrBbeRlpCWoFijUxx5W3eMxt/TkMfkffyrq+nFHKBUqgD6xB8ApOuB3/5Cce+n
j/v/3r2jzZAFFlNHGwrIxOPZD1ZXZe7pGXsGstO0m9KFF/TMw2tY5kKKlZIyN6M+3cXv0qj8NSBq
kBTbZy3kGg193stQUC21b61WMlo7QYYJ45txYCd4qze8nKjb6cMWFG0wrzXMuRWIaeFW3UHs9IB4
22tZGYGSlQWwwU3J0ZUt+jlnMVwG+ZUFZT+8M1uVC4+FeaNluS4Qv6BjyD7uQBjhL4Ne4GZ/jR7u
j/s+tI41lOqpeXofDMtqeWtbW9HxwE5Brh74FKoQEjvq2x0RosDb3rl/TSbZZA11c55ENY3lz9cx
ZMjRyQ0re1TAp7M296Kdz8gLK8qeSCTQfr8tBjar+tXp1yf5KxOkg+2+DNQIai1IAG90kcvglnYE
eeXt1mGlab0siIz8DMdasFVNn7fWwBOIRfQGubQR7BABvCgt6kKiinrxabtqazVM052uqEhsBwC1
5ZME1jsM8Z+r8SViD7GdpL10lLWTGqg4etLJW0a9Oihr+8900f9RMsbvYz7ppd3vs6Wr3J8N3Ke5
oBp5DASYRnGwsyBrCibAUqW9MaRAmjF3V/F54njpuJORGZox2djdAHi07SWYjdMCsPWd0SuX9s8T
6eJ9OXJbi7ttzj4ZuJxTcX2XhVT42OnLJF3vH6h8JC59WOMqpax4XgKP2b/4Zqg1nv4r+zGGKMaZ
kHSEqmNUXr0GI838X+24DdE50U+jHIFzWrprppw05GnxNELbJt7tHO3YQL9MamROcxXBVV7sm7UD
6B5T6yRJETGUir38c7qVuU6yHPNZCvLOOMXQVmJQfBG9S/6RcMOeD1nzvTj1NNNbgrV7OEaRjVLt
OJbsWogFnNKkGHjJVLmI1YYKrs7wrVNl4FxEuM7NYMZ8YZXfx+j35wO72X1yWNPlqSIxUruzyWHC
38rFWry19arEGxkGmq2KlQH+N37IAkLr5ehLii/8ihY16fNDMSIaw2kGYdXNeFYJfz2um69VF6yx
UiO81M60e4vaOfoZJHP/jIu+5OrLwjHZAfbM2Xcx+tN7utf3b/fTZCWEYjsgJdIJCTQ1+M+rDW52
WKDUSQgPabuGkFwig3s8QaKWFZQZkLI7KMIs9HItCq9eKpdgOjIhaBu28oPX3x2Sz28H8v3FNUbD
JW9L1VraPYcpC7xYF0RNwnvFAYQ7gLNapi0JSA7gFcEWBV1IlJAixZWd79usMRyqIK3R6/T90mzt
ufKWD8VZ5GjjRbimnz/GTKt3yBAUTITEP/HELMS6WSfOFPW6vf9wJpOqLPNO/xYQ4Qr4GeSbE8HL
EzaTr0/tm3OhLS8vmWfGLII0jzk0CG+8KBzpT7+i3lBSCy0ECD6xV+2Wo38cIQyH+jw6YrUXjJsL
cY5th5d/qDOG33MgzXjXWgHmrqRThYmEZM1TsKhAgahmahS4pPRLEyjXHo610tzAAoxBQ38/m0be
XLE22IiVzPs+inf063LFFCnCwNwUIzF+1SvD2YXvrbjkd5fFnv/4UHlW9LiZs9buGfJ4fitbkclT
IKYtAgzah0bHiGZPCY2V22DhXIhLBxfc4CM7R8cIsfcskr0exuQnMSb6R7ixReCmcSFf6M4YEPHb
MEkclSBUGtoprMWkJFQk6Jxj1NT5OWJUhRZFCF3biPySxZfCC7iW3HBLRAeH8Ins28hJsXxLjNFh
kuhGXgYSPhIexWAiw381d9Z9EnT0/VOETcLtNo3x6SnM7yT4PfluljcsHY7H9TuKZsd3jlgGT77E
bNf+q7ku7YzE7Ostkktz8UsSDwxEwrDjn1cI66MwIKoALlwMPd68TtULTXAtAHPtEkC6d3G8jsWv
ayJKBstiYIk73hgDMRm8l3f7pgKFlsuXN4Egigy2bd6+VrvvfB7i8PgNSrRg/d3SBGmZOHzV9O3A
7clKPhPG7b1rUaeM71xmmci6MevevmK4OFA7BtMJq4bZ0EAu65Ru/LcPyLgAjBzgeINUT7P0190X
KFW7FaGwaCdms7/v55x5H1mH2Zw/Jm00cq6nOfkUEeQa/riIi6ahLtRtlRYVcfMfGFkvJ7zmKnkc
7Y+fHRNt/5aqGs3t0HsRNywlrc4+9Q4sMjOH0NE5xKjfjNwicinqYY7rwtOqc6g1f98ZKluSBHeT
YYuZM/WeUCUaWfzqd+YkNjoJk7kztby/M+QzRUjlWtuvs7fYAscqs6MVQy43h6ZDBVJMbkyT5BNB
WKsJTfcZCZYeRMJ1yjZ0ouKmzbIJfL1HqDYXIfW3Er717F8abriVL7r19HCp4vETEIEv9Oh8oSQA
HcHgYVBzRtKOcfamvnvRVcBZFx+LpUCSztG69K5xksK+BNN/zWi4bsfJHaFpEX3XyUCcH7LE8E1L
3uCYMtTE5QgQRJ4TooOx6V6CRk0OFGWFEI7Y97o+y0YmzFmX1JtmUtkMzUV1+j3P83rBjAg/myXa
TqXum5oQgbdKm/cYpDA5pk7+fOtb6MV4UU6/ajjxfBcA7bvS6xnaLrL/6Vmdcg1uiDtgWWWz5QCX
KMJ02mMNTPUiq3hpRaiqFsx+p3OxCn2KW/DJnK5HyaKM7XR985dP2aYNnlROaeBb6d47Z75RmbmE
1qCElZUJlFDYgm7hQ7SdyK+iOWwUWFOv9Ex86ZORFykiUExEm/ICYV65l1XTsqQ21H47o5QJ8WQ7
TyPEXgzxgeoXCrHhZ4qDXiJlIE047yYsGkyWZDuIj13vpHvaFEXuMme0UYhYp48aWWHVfpIc8jR0
xjofjV6ykSBHDU//NjQcFs90eHWIOSVHk/QhdigI4/ufyixvPrjtwJQhld/adP6uTcbd/MYMyyDU
DwXsXr1Jqyoi3ybB+bRldo7HJ0HlH2aRb+O2NS455XCHqNZBm74jY3z0Pz4QO0hjHrkvA4Zik/bZ
D3xR+L6vbe8gcXfidVXtvbotoGAeTn+m+rZjpfClcBChHdmLoU4m+VYKRbYEHGzOoCo+iBZCs5Z1
FHzLlCcOt2e0mRM/4fQUMUnnE7QGIsQF49+Fz8jbiJdDvp4tNwOAPpiTYTJoFb0SwY6JW/4k5zOV
AOUd2neYl3HDD+1YK5cpErSn4/RQ91oG1vZepPXD5nMm6gYM24eoU8Dgq6Ivsz4X58GeVmYWzTN2
ouJG+hyRN/0zSOj8piCaINY76vgaN2pb6uNVcz0sIaYpp64+p1rAXMuxtHZcEm3pbf3saYUFWxtZ
KUIRvRw9wjNaEjFtKv1EBZUH40vqghEgbmiNLKebaiSWzCdVcILeDKs0h3LloDCWDhKdOJxtk0gr
l5VtXVEmamb+MQpCA+cPsM7CNsKjLs2kN8dN5tyWXis9TrUB4v4TKHIKTjOhCd7ARDGmRnfeWMwM
DaNFHZPhEqwyDUut0ml6gwSF1A+/RVRGf8GkZyKwD65w1oj8jySe6ecPthvXZazmlKHnaiI3MUQO
xfsZVkVD7t1yzDDtauMJ3YOjTq+Cvkf6okfOkes3rZ3kJH8azqOJY6tJ8M7B+CJL72+7CJcJYAhI
LRzlp21Echyu0HFNGAaST8oldOzIDMtk6Z2NOvg8S3GJCrV8cycXrH7Ug6QbOQgCf4kV6cofGwp0
1yAvi2IVoBW5U8yo3u3bTgukJqxVePwaOYkppcEozNR7zjsRtHIP0TsJWbiNNrfKHOOBKzvrnXwZ
NpUU29WW1u1LM99D03Ypm4RxpI7pF5z8AToceK5hx5cdt30I1uEC+xiAv2cdkKh6jzUfkqWyJgWZ
xOd1BFY8tjcyUpyapmZtm57oDSyud5xnuAZb8mPRj4xuz4UIxQOG0w7O9DwyU07gNtvr+KWL5+Sq
a8biuRzu60NGVSUosgUxM5cXQq4ZNXxCYesf0WGmrCSouqjI13SghEZUCqSqbV7QuUqhYuO2P2Rh
1YD5/QFZanJLejstFId3WHyBbOOyj1qPN0Iu72uFYXvA342q67b6BOw87wcUZh0Wi+kgGVIfFyLC
AHrfOauRrwFOkbNk5AB6mf73O9P5/ck6puTv7s4blQPIUXxoJ9iXR4mvdyPN8s00Al/kqyQ+VRLg
4II4Fr8Fwryr5dKo7O9bXiwMBYqlz7cxdurBkk8XiarA9yl42A+l8+aBhI/940sL3BcfLvccSNAb
v/Y3PV8ydZbt3KSoBQLgndHu9QE9kaQEt7YBPv4GFJ3Qk5kxheIKNqWKSApixu9wFCF/jL2weHrv
Eig/Cm0dwL48u+a8rvs9z4Gff936NtWqqm3+GnpTTl+HxaYOWwStKvJKRH4KxTSa8hL1VL2ZWYN5
Hyd/yRL7+eJrGB9dQVvtpmcemVJkZzNGM2T69uLZjQ0TlVh1GHC6D8XNABbkjXcKTL09Rr+B7tT6
YGtAYgR/TVW+q/g8H2yYhed0ht3pbp5WYE34w8GtOVQ8Il6/IDRYgU2pXUQ9xbVUMp1LhWnVpLRT
MHaRgZiQNwV9xtIKwJ4nntOn+KxJbcb2V3Vw0lxzHoPD8jYmz/JwRX/QEKb0Dc7+6H0eKgdTV2Jx
Te7As3Wt0g/r9AC4LwNynDCwjgV14kgF+OxLgPOUh7XCFz3LljPYoZ7YYv95mh4td9WVudS/yWtN
vIeuREgs4aWmcMcE5p1j84xAqSr56nIkc+7pZTXiLOmDb35JUc7f9+HNglahPFlfU2wLaXzJT5UE
ENex1p1Ya5QYT8xoJz/K95l6UzbIq8k2GK4q/zEWALHb5IYOQbDVys0ma/YbH1lOf+4P0cmrfSp4
2M8cPiGmcrE7Jq9azI8yW7JySiLOcPkXAXK10mGQvGxx4ZaR0DN1zyJwhuZtYlqaz45/RsDoDtNa
ik94F4pMOhfJYISI+TbfAjMspeCuK7oIM8CIVAXhVFUJwAim5lgGrauCsGSgzlTCnxJu8twL1tH3
LYsbn7x36HhoBFpZ5/QzVpi8/LPDflS1O8+UU5BqGLgFp/HLxqKp5Ct62O4BySwECGM/D+7aCbho
INI1TbPIuFoUX3XKzJAgv3upVUxqqvN21lk99asp48OprcjtdGFw6owhpWlp7PmKVlaQ6dvR8PVH
MlaYNLTfbFlmvLSFJPHFlrhVbQwNh8KiaV2T5XMCD4kgltCHhOgX1FoQf0sCl2h3RH9Az7YeseFv
GZ/C5kzTcsIqmV4pmh7DG7v8EsSHRrofeg42hpXtth4Ddw9S9JnJtfnc2KNREVcsNXnbDAGeq2fv
D3/La5Go70PUqEZEe9baFcd/GZ9E+u0+aA7Gvm1otoY58jvGFrbLZcChq0CY4CYV3Uh2xmmFmBW5
zIN/Ov4/dZMpATeW+0TIex+ghuAw+ptyxAIkgqU1GdwWuEXc/yGPgJ0LM19nSNfYinvWh5Vb0dQY
ShhynUsmza/WyfHbBRCqiiuhqab2pQpk8X08RHYkf5p67Q0Tv3VJvzyFQglC7wLUJMKaY5Fmtd6u
I397VlN9pGeAPnrDPD3+Tb+geNbqI7RGQ+wML6Bs3o/wR+MnQkVFtMfTVuY5FXPZWRJGLhkNYBGo
RGulX2LhvcRQXvNyYruVxAElVHElNTFGfPz0a9CgQBb/PRnmC9Skep0awcGZbVBOwQXsCh18Fvk9
50PPQ8XYeAkGPielL557eGL+GpRgFhh3NTXQc78/J+J9M+d3Q8NWcRlRlDOSKgQjv7z9H2o5QuYB
QwelXTn30kOzBBNRL3T8NX2XNZ5kS0mHnLHuiFK6V8SSujtf40zvjBMK46BFbchvC82l1gHhvN0B
H9QqBOur23jntxlHixZSn4tGrh2szG+wXwDkpKbngsgPOgFj6Av0TN/RTAMOo1sGkYCbG6kqcC78
8qC/hDjXE7oN6vbTOEWFtJB2zAKnduXbe4/c2ldXYX8SzH7SGpIlC4d90QjeEHxNLo5Tr1JnMwk/
tXo0gtC/vqQIQoiXYI2ri2HHZQeBSXd09+8y/Et7Vnyx58CIYRTYi4/4jQgtDpfMG0nW/xLZumUi
IT0I7qT3fqq0WBmR9VNSJwMKcfuuHYPEl6ww2lTG9SXO/cCCl38yBprdBlDRVTaSXUUwjc8/nmrq
D+A2FpLMUFADCrYoex97lnVanPSrCsK9dnLqU/TkmlKvPIanJlEK4m+7FKIPOtHP+PR6PV0a+nLC
wIWDQSeuq9Ealc2YiGlDavoEMmfPRnSOMy0uIiEa8tRhz4cz5VIHNv9s3yfFxyvyTPjA+5uWKSBv
fgn4JNx9HYsIcHsFR6rVm2vt6XmVxWAR42Kzwddp886qgiomPlShmlpToUHNno541oi3qPS4yRWi
kd/3AEPVafTsbHH400sm+9axa4aWxQsKxpQMDGrGU64wmLar11wAvTZs2y0jQuvgpzexzRsGiw6H
qZfykYj585o3c12JFmfzK8Urqvm4+rDQpZyTZtKqjA5sq1bpKsQeZs75ZBOW19Iar+SG4qiuy9Ka
562eZLzFyuMcigVLOPKLxiBU817np8grfOMA8ZXNG41wVtUHJLUZ0AF/ndNc4q9bl6cq1BWoFv9Q
tmgj7CB3+MYXryYW30dwNPnaibvOx6sOqgD8RIj1Lu07XXSkqITaGw8Uxotmr5mXdaifAboF2YvO
ytP40Ca+RnMIFYGyFX2oSnUsWFPGhrdOTrt15RiVllE17yUJQSgy+lI2Uv7svx9A2Am1sef5o/xV
90wdq7JwooSaumHjwOy1AohTNhX20oWMlHm4N22PIUgzVy1XUZtIJ7adefkJFQlNrnKIK1wcS9U6
zQHTEeVZ2CCcJ2FIGWXkE9lDIYvDHY84NZ/nVRIH2/jb0SHB7XcrfjA8TxsWO2qQN5cUhKkNWlZc
9H4hUtCY9hOdyqcLXzhWshIMvxIOaK+gc0WIhqu/BBYfOZU7TILk6XdpchHgo6C0ejh6vnhdZW5N
7XyEWWzK4IFx3A+89J68HBq18wKcnVhaLgScTfuhCgNSNK7dTdzKXLmvaHZkD5eayhQzpn2JaDpQ
VB1fZdBPSeTLZsfSnZ1ZnY8UZOkjQC5zVUZV5pIV/EKFBACpPkRUkJMUAKMi9mPA0cnKbaRACf+9
9hWVji0Ko5ew45o039smsd68ChjrNf9vVYRlmLF8SY1KoAaWgTaEUkvn8Jl3AklLIyoYZ3xl0deE
pWI2IOUBD9NjAs4tMKoFRD+b4HESZwnidRkU9pKDXRtEMdlQJZCrGdzTs/0odiH2mQyWVCKwCWXn
QWVHwSWlXyfc3VmV05+1Xoiy0SxkbS5lKUvTEyHS1tpcQWmWYnhRqziZLO14J2HxBaYVPMEXRIrt
o/kUbjrs38ddXPkhRk2WhO1WSr50rP3sw6lsSV34ZcBFyrY+/4ebrke7MY/++IWEJOxpDXbDiX2M
3GNR6pBFn5gio2vvBBIr/+Z4TfpI+QEVN59CnZ0sqBycqhBfJ14vk2j50D0gh1scPBURawBrr8UZ
EQD93rIiJRyFwDqYNWn/TF3LH8m37cGysXmsiiH2O25WRPFkbR8qdtXPWUOKwC7T4rHw/QO6RL0R
6OYUzlv9wIgJxDDEqd7/4fqpP0REMejnBArrDiyFQzdNxsjLI0ls2B/cNktyDt4MLBZv4I8tmZt6
ha8p9spdePsHxNCGg7+PDwdjoRXK0ZtfQ97WEBTXOjHR8LXKMhaheOIq6cX+V3qde9jdHbaPsU9D
WjHWNgq7P/AiNX761Y2CrMPeB/uz1Zp44zUsn0jwF9de96baftyW/BV13IRtUuq8rsf1MuGusM+y
z7z5rgMJ7WRZ9rQqTZfoBz4OFgtScCRNuYOEIcc6uYhjkLRl1u7rPStCxosEoVuZprUXE6tsYbGj
AEKb7/Vug67jZC+wLZhnLgffMcf2d/kTOHTpM9napOdTBTZpTGNkdv//bXYxhiJ1/RQRrjvhRqPv
XNVdPEsAEA/mkYAlcjt6u4xst6vusqNJvNrQ0ea3/1c7mhjXnjih7ItEfEmloTji3gBBrt4BGGki
kW9LnlVmZbj1v32IXv5sJ7QY9nN3+iGjkDFN9xn9P/PmhYs2pfZZbLcTj6lFyX7/HkH1W6plEFg8
tZJ2sKMJwXgqbd5qnoL0hfAGreMck+lG1bY5dSfKOi0eX6voCcW2on+kPh35byLE82u2Qh4Kbf5I
J0AeTmsWM0nOq/AAs0POJvSCl9Qmq2htGSnXzd4Bxirmo5xuzw7J+3F5wJJg2nJnzHp3tGVL+uzM
meDM+xq4ok1BaRJFWTKF0FW3ZvxEAqyYRsleVCJyKMprkuAIrXrmtMI5duzx2ld659n4hnjk7THL
emOxks9OQl92cywjrDHld396ev2ivIFreUIIxgaFf9fLPtwYofeCVme7dXcdfpVjrHa/rWjfJ1qc
uoLUjJ7MBnzfsStAk+8NsQwK5FwsCWPlJ8Os3YIKxxVV0yZGesOelM7rXFPryWrks7AS1TVgcxYI
g4A4BpIs4ubQcrG7Ete5574PnxnkGhSF47cQ5H3eG43UvtjHWJnD9AfP/5N5ftx0W/F+Y9+VadN2
6YHd4HpSC0KKoiWUoe2xFd7l5O+sKaS+1mzagaDspzNCROOOmb2H8PQ2kcstCgxgDPImUKtL7wbP
AwuUGZCscnKj42VqZIl3ZZidT/mn13eCc0PurI9IfBbxebXVtV/eXzF+OQSjwv9c5YDhjrsMKuJS
2YT8gXbEWlE320y0ZO0PA+v6iuh4S6XcuRA2YNprlQUzmv7T0dK3SycAcBe88pLQYy8UcpJWI2uF
5LewTr/37Mz7lXWjavlUCEvhuvVxNFUB749nBrkpU1n+67vT9qfJjhSTihB6yxvAk3dYhF+uXaeE
Q7KIMVd2Wy8K/QbLHsKipEi/Dw824hH78X21CZ2xavovhLLYQqnLq+WF4hsFogpopZ3FJGjY5zFN
Kci8CTRXeLqVLLduRrcNzTiiZpdmtCXVuW3qKkC5q/zxw95KJ/Tz/TK3exIjli1zOrAgfN9rh54e
TjWYlwqUJfAZzHkxUFSCbW3/MTfVs8UCxnaVPBfe3vqOQ9ajku5pcQ9nqih2JkCWIEKedkbjxB7R
XDc4zWiJ8211wM2hkzlpXm9kSzpzbonIEFiBRkJZQ8aJg8pR3LSCx6HrBtsl7SYgaJtyaOiQm1zn
1xdjzUJi0FTE75ekYSBkfvyEsTkXboypp6/NPmIMuEujwCAxYdZiQB/7fHfKyMQISKwtsdhnRFbl
Sg3DTXEqHXPJPLhGJF/brOK5k/ZR70PHtSEbp84VwT1MxhiOteQVnMXL5/xDrj57oOQ/WuBdI+eR
OOWVLkTz9JxtTWhTrEr1j9X/cZhc47enKL3VAJWTD4ZP2NO504HsbHwAthEmudryT2qamYXPW+8V
GH/EEwTRaV60CADLeZYao1Nlo8Nb/DY4Sa65dn7xttv1evJhgqmncRM0xz87a0jtagaifgKSdtbW
JVDsUeZ4yZLSOnjZ8ZVoLZXawjZv3U11IVLLpYGUN0bUZw1TcnsuDG/30FD8EZinDs84RdLMq4gD
B/xxkON6DRJ3MNePN2D66ePXwTOWO/Eg0GD8JSPvZX43rWLyOr2HUlHJFmnq27V0N32Ruts8VvT3
+mPYPNLShyOnVW9T0wbyJ8SCkNjTsBGN+/Dx+3B2rWu+HtNBs29GHTirGatxXKpTF3IYDb/ABYeQ
qYoUi7jB5MLBFSDN3B7cTyG8usVdYB0St2W8Fngwg7xusLaKUng0sAZIbl9sQ16irbVC9vjGjT7q
wCrQaNbXigX9WxYB4vrt0C7y0cK9jCYJj07hIx1e+L6U+mQ1TxCioQ3Td0AP5N49CJqYCXDqYxxJ
mHLyTF0Q2OaMFTmBbYNBnA4qMUopyoeYt5daAB6TVyMkNBNdXnX6McZmQqxGJ0DBXzos4GiNVI68
Th+zs8frA7ArI4mMAOtRhkQhGOFGLHzwLxPLP6hsX6ufaDHr+kKfM6E3m0fQFocM3gVxyvCmdL57
rbT191KtQGDvFkZv5juUMnpiu18B9XKN44j0WpHyPWeJEakaz16wfzNoo7zrqdrB4yMB4VFTeYFb
eHzTO/m719TBIB3xOOFMv9mS9sIBJpM5/6KsoTbKLcT0z+jejUqdPuTPcxdf2x7ELsOuSdBewwNC
lZm4TpBHCHtqwC071RwPPjueBF4BQxFajrspskPwhoAx7GGC8xASiehvoilv0q4NsAGidngI7Frg
Gc26wl+TwTOCFdw/aw0Xs/Ey33YlCVmYh1P0vpofvsGhu+5ee1rQUUkAGbSaW9PMWkd51FmbJdSf
0W80FUXb/X6Wb3OQ3yCs6bVUQ7eglgvFCxwU7hhgCbQ6jxln06PQyNVJW6W4h8L2ja7j6/QtzV6Q
uUFyV+c3AOObuKyDT8UCWDNHC+Oeu3TMjtj1D96os16wzF7kqi/rJzMKE9muOmioKntuWITOrq3X
c6jHd/759Fndrfm94F2nXMbIN0Fpa6kx65tNk3rQzLyRmISB/p6jPyV1XuejGcmRFbCRxMXYWMxW
em6Yh8e/hIHGLqXvOp0/zM+jrasclpv9GzIP2RKfmDePAJ1acfqBpKRQuMz0jdkyr8uPN9J00AKi
phINE2Fz5D6O/S0ie9QXNNpSIvfK05JE3e23ZfmuN5MDMaQpU/pxmc0PN4jkFYz0uAnoTLWL4Uej
j/qabrbMprvnG4hO3Rry2Z86JPxcfUA3gt4cfby5CXRo2jricg+twITya2lJ7/IobNsMhAmU/cD7
vanTUJrfLl3WMbRTvsOMKU2Jc7mQdCArtv0ShoS0r9MwUZm77LUnrPgcj2RvqSiCDna51GljcFE3
EBNfDjh7WjHSFVGIykEdluJyhsct/3jUn4a9gugXErG/zLZwaXGA/y5YJ5IgOy5iwXPO1JwO9YO4
o445totZfz/ewvzYmHzJRPAcADwbDQVXer8hnLTKFkKgzKDSTYQcWmC4hQA1NEwIv//4xQkgWmUE
crhH3YpOGAaXLERA4SNZNjZ3A+ralpXock0+G0cSQT1Y9gbBoRzhzqWdnb+ucjbGVOQueWGTJYIx
fR3rrzEeLcH9KWGOxUEFvdI8DU1QNyrw9wVYHYbCx8OwFuENLZz5gVkAHq7Y47BYql7EDjO7HzjO
Kvb7rY+O/cWmFE8jlUXmt3YPrNGCWUkFhYAIYWsdGuExB7TcrUY+tsatk/zZZEKLIV8YdKFewP5p
KxGNuaYwe78hs5/eMm94WD+hKQCM6V8G7UdU6Bu0z1MEDiFdaQSWee7eD03BnpLMV9zr74R5yIrv
X7bZL1WphvkoJGP1ntz2GUW4z6jHAlHq1j3wGzs1i2435n1R+2arGhhzW5+tiBIvmtARVnXJjyfl
14oODrSQlafu3GMH4tlCKnCPIbt4FOy70fC63C6YTYIFALljIdIKfhSF1P1NWJHIe7z8wglafekK
1z97mOja7AanmVbJ20F8buz/l3g73sRe7cu1+8uVZ2VCLKJFFVKaf3XspvMNkPt9LQ4I7zylp7PG
+I4sHaFxi3qOtMLC10LhKXPy9ZwwK/D2MqUauogTD3GLE/jT7hEIsq7P5dOXPKGrpZu9T2V1U5/d
RzMv0X2KladZVBtS2ohT3fbvCepEVZZZqVw3MCGIUnPivnm10Q5nCdewDjpW+N+VX+yU0gO8Dhvl
FFYcyDV4BOPYg8JJ+iySrks1pz992a4nqLWTgBECi0Z/RUP8PYMwjGe2jWcAdWgXJFviOP+Q32tI
AIjhj6j7rSDDL2SusZX/hR5K3oxqynhudkVW0kYDV6iAhkDXe6xac6FwOA5k/qbN+22y/h3sx/ZO
gcWIJHj7tnRefR4bMv1OGUsOSb0s3iPmCg+68/9ulFYNACVvFeR36LexAVvz2NEiu6WG7pHzgqa+
+4Yw09IWot1wxBNowS4UoXdGRh49wvZEowhRIkwS0Sm52uDMtgR3F1Umb7rECmudoJ9E4oYLLmCQ
tyPWJ97PzfIW0PQFhYjw6+F2oPfNUU/4HAtZ3zFUroWFeRpf0Kd7RB5pX1LX5jXStKRv2G29Q+/w
JxV4oQEQZ7HSXENmwymh7qKHh0UoWjjbfpapjYPAna5UDnehwGMKHDSLNNyFfNH9Qcbx4UAA33x8
cCQYEkHs6e0PiUR83Mz26e5u74NGkwCtlk5EmrW9UwuBoxmEALyLbRxE455OKDA/lTVdHt32cPUr
cNq5Jgg20puNhcYcW/ZtITMxJulTOp2rYaBXuPw6DyeOY9sWxlLK94TycJ0EY62wc6ycD2z7oqQn
sa0iQJBJ5ylijATx0KgIWi58seWv8hG1c6QXNcKHCcnGsjTejkD29LqUUesD3VZkj1clJjTPN1Oa
oJBFkE/Zz/vbRWDof3deQxDysYQmh5NUtoRzbqZP+qkbxMm7cYtpZ5Wfx7ZzWFNMK5PKURRfUUoB
UsBCFXB7D9I1anXgsZYC2at9a8EiIDIr/wnp4Ck8e+cCJTkDwrqs/nBAB8hCUtk8LmlDe3gz0i4v
Y77fCj/b9NvvWxLM8Q2Jmc14T8XdHkzYyL3xiG07JFp1Zm7u165RK9UhsYVENyER4Rxif0IFq1Lp
0215mbmWp+SbyUs/3s/YCIS0Q6Lutb0itkzon9wvnyh0qmjpkB5vs/9+7eHnwSEnEdghlyJIrTs7
WOHaWB63kVzJRc2/mrVdBadHqxErxmmHDLzlQQ+y8N3iX5WJNH3e/CKdAX7E7ymcn77C63Jfkspc
0JBVKw2Qw1QJtzKjHD4CE2tFIvY45wwqS1xPGfNrG/zKhst302lQj+CdID6W/H2Hdixh2tgQP6g3
YnyDqmSiqMmYxjydq9Y5FMZpWx7Dal+1ZKRE78nyjn/ZY/u7wl62l/FlHIEguSrc7QnLPxSTsb1k
JC2OBeXylqC312DVRopYF8QsOQePtTqtQHrWmxSgrK7Voer2R0VcRe36508VV+4qpsFFpFOxwhAg
IacHi8GhZg/i/5uAhL1Lgo3CMs/o5A2BZspckqluxhShJROmhJ4Ln2Xa+ZLERJhwO2kWMZZqv65W
FYsKR59GFxLc9MAEEq78S6BxzrE4X5hAhfdClkoxaCbZD2Ggf6zs6ZcKizClXT5CITmIwIDXe6cU
4uw6nnEvYioRnl9P9tbKLnmuE7VmtIms2rdV0tzFxCavjyxzkSsXIlS+VQ6QFplUGWEPDzg4DKmP
dUl677vTv36HLYPp5NA0VkZrbIzc8gTdWe96f2m48WzX916rbXtfxYk5ibYgsFIgIWNsNsiyGQCt
xzqiM5iSaHzi/aJez8R5O1ECGe/6jV4sdy5tL+DczHITLHKAans7fhhuY/PodwHQ42GBkPk3lNHT
z+7tg2otevdFUnKOrwELOWUbQz98BJVkTWgWwkmKRFQ5oz+xuxy4fECBWCTJNbbrc2ErME3+9748
RXDJwL9IVK3Sha51usTAAV7U2LUO2Cg7aEw77blcJotsuG1g8dgoemPgJgUsyK5e+2PR+ePF3MMy
IULsKnN3E2sE03g1A1DjXUFByI8ul++oceqTzZV1tf8kT/7Je1Y4eflQ149mWL/1NRtOBVScoJPd
LKXYw7K4YfTl7VlfvhNwJ16QVzvjd94D7BmqOSCfJh1dl7TclUJQjoN/WNvTxhsuqqbdEKau704c
HzegHmnRvtE1vulSY39a5g3T27ZaxBSRJFMR3fcHXrsfhQ+k+Y7+JZ3wuwAYqNwLed/HStLahEQN
sZvtbVnkyuiG3iCIkcRWcj6uliaCLcf8nCZTWOx/bLVXhDMktpO06ZuMo2M2g18WGFGCSHB873ua
iTUgWJGueMP8ozhuULWhV6IJZ+J94GxQgHX+knPvB01QlqDTSW9oawtSZk32R+HeFLZK3baCnYiR
psoAkiIQUGLFQaXiAskfoI6S+m9ttDC0eYb+cJ0MPq5RwqZood7qpJ7PTizuE4taawvV3aHoXq3q
GMHWvWVKiLeJ5YSYJhe/lThB6HrRvvPTuCz2Gn0P1P0QGA1zEeJAM6FdAaDiUwRiVbCbgSMPPX55
TgFmvS4vPiNtW0yPPGxiAgr8YbUnnXbdQUn3tdmVM9fBgVH11c9YXtmPcI32G9P1HW3sLMh11kHw
uJuFBg7cUJEzgM6FjMVeMSd162rzuglU6JpTdiP8yrdGZ+xAeUUBaCkl1fs0V9ex3iwFsAZWSkh0
zcnvRxBxpJwhBTX8M8IR+6ZqkgqQXIlejtO4HIHydjIcHFUqvFjkyidZtKPJbIyirn0IhBy/pZHw
yuVPdA+cj9yGNs5WDZ41Tg2ss0aKm2ykJ6j3YUHGOdX7p5ZCim78EJeIiUiFVVbldxAfeVKpnN7b
Qdm8PM99Gil7Ix4ILbH2j8Z1x91QQORaR4U56Hr103BXvLgtLEqak72hRPPhqgxzWGXydu4lonDd
cqfYF+jYuD/Gel2b+KJN4Oj7yNaTwHUxOG/weMMH9d26P7w6DquHxf7l8RS2eT4KmyYLgGqt6pDW
W1msdKWb0hcx/HOGTkyy24hFlUZqZJSuTjKhsOG45Z1I1nIjExIeuU93Kp9q8oYkl/8ZXD5BRpTG
f2kdY38bp/JOTdgCLVAVKx4LXIkXcQ2Hm3bH/BdWUL8VBQZawy1zb1h2d2ipy3k2V5mDel79uRMw
HTB6uqr0pPOG2UqtulwWVFrPLQkPZ6vUWlSf7suDBm1xq60rI41kdJRrCbuQBPsYXS8UrEtR2kzC
ZorLG7ZXVxqIGzCgtCI2mEM2ybXtl3P99jeVCzXrZiDH47dlGK2qi2f2j+d85evRD0icgty7uyPF
DPnF+uCsJESQCk7gj8H+Cah8hm8Fj9hU3vDJf9eH78Z4IAmHuRUgCw4XVf2KXx9jOtUWKK20xhCw
UFPDrEcUiHdCgtOWT17fIBq0kz8/55z/BEnM3Jsp9c754o0wKl7iels6MkB0tfQdLuP9Xbnlbj0b
Dme6m00ItnjjdXJu8KtGiR4+P3n/Il5f/8BFIGW4oQEhbsoW5Cz3kc36UC5DGETnYkP9mfHOboUt
OPf6gbWV2DNTCWVsmH3Yx4HluWifXwQHLftknCm3EmUgjKdRlnfCMYC8cRMSkTcXrmBErA8b7UK3
4u2PK/Rc+t2nh/CSS6WzYsxFxVl01QwcqZC95gvQDt5dMf7RlhYjt97cKg4P5opZ1M5OFE9BRq5D
+8UkuUPgc2RdgoWZk/YSgxDeYiFtyrqeXW5q8e0LDLHClYNGtO3cU3SG8euGeMBncSov28zxtPwv
F2W2AtCSTmMv2R2FZgGOWrGlDZatKeKYWvifk1nmTHt7cwQKM+/3QkfisyIdQwcvxiw9lgGlj1HB
oLHJI2dzXSxZNSposvipqJWzKf7ZqCgY7k+qVPoqqDPUcVgEM+YpZekcOMHaG29xOnMIKhCikVDI
YV5DeEgS/og9kQwWJ3QSJBhYq5Yzc6BmcJZP5K61+Tx1ZFHoIORuz+PqNDAO2iJGHIBaC2quqDpC
cloT6ssgVgVUvZutlnLc8WHXWRhH6TII/5A4nv072uRR2qDZ6+iszLkVqGUl1zJHfupuOQKZrMqv
TFG5JxOEJokL/HXJucn9Sa+NY2acfnLB8oA48RvwUtA6RY6fQO3HjXgjau0cy6XwKVV2SN9yGHQT
3ecKrv3EFK4fMbaAz4+taz3F62/6dTCqt+WpojqJ3BSOEmNjPTbpR4nxusP3ZnDa2jvq9sTN91TZ
50ROMEaMCSbR3JEKYcGERLvnAx7bBVJuk1j2MCuBHQA8PDEw7KhTUc+b2isEULymSw0RgKAIS+/u
mrJeqdzcv3qscdkqoW4vQQDnoSmUfqtRIYUhszQtXhwy+NmY7SbtDp+YGbUggw1p4+NZt5oS7wHA
94cYF9e8PjqnNxhWc17YxCVvloye3VN1PJRFuH2XZypT2D7rkiR3irjJTfLJIrhY3nXnpbuo00tW
uURAVK8Ci7Rdw367sgO3gPbMGE++9WjRLYkVhAMNt55GTYhJ92q+V8bpvBtFzIFAd1QUPSY/Qiix
H1dpSTk9ubtbP3Fpgutu6aRrn+PT/cutjtuW7fsAi1gK6cHcrag21z9/W/bFFEgb1oLs9/funE43
3GzXqG2TrfehKu6Mz++5lakHO0n/VZJ4Yj4jvNnb3YpK2Hbp5ebrhsXvzS3vIfFEFBxiVIPajTHd
b9s2tF1JsP7ebJICtdov3QMAh1VExgXlcC0aqbOuGbQBtqFmjHV3cie7vzq5/UvZoc4ZC1RP60Am
f3AIRUACG1gxITlZSdk0+6ct3WLvilPm93lgZpbg3fiQpZFuVGatQCFBPBL7/JeoKf+UOyletajn
pkyaNTzmSgCNMbHBFNByLIceCW3ASX/O9qLNKaTNPlLdH81YK0ldxSJ6+wXtGmJr8sR3cZb04d+5
mUs8CXE2mAIuyMX/hb2haIyT21LSnURqjscECakJ6o3liR1Yxh038WXCBjkjGM0pXepK7kEvZYPo
lynvclMAsuwJ3dR/5FSo+lImnj2Ahvndduog0b76TNb4nCmZmSznwOK3idkm6C3ZEuwtqhtUsukm
WX66xhVAEbDZypms2Z6VqhR84zRy3UMi5FnnSEWz0QALmsDkyLdi9K4skr12uflwS9C+7DGvLERM
mU+fQNmeLZDyzpXLK9yTDGLdtMtJUdl8ywtLeF1LJ+cRw0qeSKOBy147IROVBeFv4eBa6dnjAhRs
ZgsssY/gzXKvJJkkgZjd4YHkf1UMlAZ+4BCIs2QT+ubHMmacxQRYr7KoNigL/AJSUoTqdzAsrIPp
tzNGhuCqJIya3dgUk2rSNB43PVAn7Mx8Io+CcofsPekEt/FdadzzpVFmwSSOUjydryYjjc7Xd19W
WA9bN92JtFXwJUFI+zDooRLagc513AE1Wf/Qfmyf4linH4Ur+2KoN9iCJnG6ozxe4EW/YZ+TaRnG
0ICK4w1gZ4ksuvKbFd/takZV73VvCT1WKNuMG+8Egfdxf650l99Ei+Bx8yrXPijdQaRehxBNKzWf
gdL88zuer8hII4F0N8Cm6elSBA/oOa/5kwJNa411ryj1HvmvhshCtj9ePl0Oob1g/GN2bfgyHXo1
ynwsInOIkyvvLIlsNqQ6if12J3wt3qHfqPHDJxt2O0qnw/FNelrXvWWdUuIVWNLKJkeXJ+H2Gxp1
90zIJhpBG2m8X0iOr0NoSUaFMT677Xxz1RUYPWfUYFXqMJeQCWYufF6DRrOoCyNbNB3fU5xFHReJ
9UWuD6VbumfpWqLAXRis+/4R2x+RVWU/KRn096WUF7OGxX4l52J6NwGBI/Hpt4Ad8gs91g/XCQcg
E/NFlR/zexLTGZlOpqfywOXhWav3AJvTluIYguoEF/HqmnILAcftDNXV3b3pP3KssmjU/NrgKWbC
w++NqIbXsiGO3UWSMyx953VRuN8G6RimgV6zzNcHHapK29M2TZI2Sm4bUAOWzuryzeRgrRYkJa4e
7FHuE21GW0uS/jN/6zkPnTi9TO9sWldcN9ml2tC76iQ9a8Dr4r3OcKnZh8l5DtbYQJkRmy2sDehn
3PE6X49GXLSXim7E2K3ysY0tMEBJC6seyUeIUr7lbPTIg3Dy01PSuGuRKY3s+k5CFsnCTaNBdPh5
kq43p43guXJfdATgNk6ZSmuxXLEB5W0ggCSlLK37oczr9/iI1aWMZb5sMVWD/dfY2DxaoWcuz+HV
Yxgpi2PSQCCQrVCw9HBengEooo+MsxCKqpqB4B60CfzT84ocaK2yaG3iWx5BvZo6L3ZHBLbZYX+e
q102Fex+OlBQIkZiZWx2mGamm3y2ObgW42LozGS0lufTDlsffpyW6AcRrCsbZbT0U/V7UOz6R3IG
Esl58Elu2OU1CQ99pahl+O177HPS4ELQbBhgiQmmDhbWx+rf4+gApoz4i80Veo1JcUnbTXQ0vDpA
Y9hOAP5hKlq8cKulxMwRGhK8V6pH/obPPBwf8WHmY/cyUu1IMhysmSQwWjvYBvw8tZmBK8Chhy6G
tjHO/MGhrruj9jh1/57GGp8s/9i22Zj8RiTY9ACqKvFmQiWz9zlIkwQydm8wgQ/SLO0G0B8MNW3q
xJcXxPYTHJ3hr8wqUEH7eDKz01vo/xLKNHQPbKdDsgtbNivVBi3MNTmVg15WfcC3k+xPBOHb811j
JTrEB3jProyEQXJbB74KVuDxMVv6Sh/ImcM5HAbKz5EgtaWiNU+eETaMHGIOMzQxRlIb0pQ4rvKc
oGQMWjz/Tuh8Dx3uWngc18Unc/EILYCq5vobVkW7wJuDybracq6IU1C01kH7uNt2LWUJUW2h7fqP
Txze4k5mPRBAbIzQ3hzhWdjxD7eUNIdUlIN2cf+QKJLYCQMxupLZJAG3HFxr0z6fmblGmckbkach
xroofqKTvuaAaA==
`protect end_protected
