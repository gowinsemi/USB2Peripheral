`protect begin_protected
`protect version="2.1"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2021-10",key_method="rsa"
`protect key_block
iw48CaFRpTZ+2yCrTV3WRDGPEKgXZscdORaHPi41F8sTb2+Hn1aKo32uVbx4V3BBPuAgWps+r3z6
76QTzPTql0WasJP0YarvqKYpimDnj4cj7c8kVIn8j8USxGd5OFADWFxUigtMM0miSXsmV86DK0+d
lnElU4qnXa/1IeSX9jao388X0aOzRwJTymdOW1kH8cdKSqSVPErdVIYfkNu2bmJ5METZ8RLhllLU
qEC3Z1tPoiLdBALVPMhENvF8qOqbPRB7+ANF/c6FobP4Aec4YJ0wETNc3p/YLHtf0VMXNVQN1Wb3
AE1kh9bg7pS4V5/RlADsLvP/UVMQeU8OU/NuAQ==

`protect encoding=(enctype="base64", line_length=76, bytes=20432)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
nRZLvG29VehPJyd6u7ommhF/AkVoIP3OBqCFLnpJq9wcwr8K1I+NV8ayYO4KwaVEGVl1FzQDR9qz
/lXNKwuUG0AyCjddPSqBsdtlMP0CXWlWnxy5bQmSQEKPRUc2zrCYz8WWVP3jBklf5LD+qKQq2CG0
S47uVYVzP10z0r0lg9VM1e1sjQmeJZVmGjJbucjxs2yZ+NR39q1ownTalAsC9wpsNvOVCobmZcpK
XlPXRtv5iXEDXbhW0gWTgvmOwcNZhVkWLgviyrb3B7K+hySQT8/Cz3f5957xTS1w+nkitT5JztW0
4GCXOgUrpaZQP90Q2iRdB0OFgZ8UKAgv0Jo5BNWLjSau+T9qu6dqYEEzpQmuYJJWVKSg1pK22Rwq
1F7plIOalvcyZja0mTTRQDSG0MlgSQMj2HKG4LBlTUBf+FtaEBr8YV+BtAwU0Tbj+uu5Rnw/WVV/
Tq4dURT0xCkau7T6nDDYXsDec493cIlF0wv44sqhHBY5BErPkA9KgpOSmkbOmi4qQe0+b0SmElJn
6g1TCbmCAISTMvPeV6lOAJc6fRpvjuEnqtBPyH99r+l5AQZhXqcmHr6OtLfronOBRWRcn6AKJHtn
vnEnMx5TIZPCbSwe0K9QFkX4efmbxUdo0fY+f19LWXyB+zJ0idIMy0daNQQAAjZ/1k+yicVtKotT
aRa9OBvskani6xDeM7olM0hudgIF8eZnlZ80dO+MLtK+ZkDBjV/OMIa5j+JBtBl6VYpdVHj6M2ts
fEHdc+5u1mqwBrtc01kBvkYqU7LGzjCLrzBotrLX+aqreyPkSv6HSu0w0HyKSdKDMPV4C98fZ9kP
AvtSyOsAK3szcKgm4JcRCyATrvcQ5Xu9gNbD7T2F+VN2qDNvOev6iGgaUxeJBo1HSrNGSP2BUgkp
8p951kr6yy0khmMlohlezxTt+5I/rRiV9pwTBxhe9/Q1xy4GtMc+81aT/qckJq0khETNcjNOtGnu
3mIT1Pz1Wc7Fc6LyiVHhE9yw3hI43jL9VJBf9O232yH2N5CuT6MbZ4Mo0qgk0esMvw69foDIPEI4
9hILLS121JttANql74i+DU4h5uccY/7yZ7kEGDV5wRu/tUWEJ1aLe9gpSLeABuvYHzRyDrxb1HEO
EkTBEm1zSlDPsGsCJKs9Vc3kIjKNCg+OHcI6WoLNke8DVHvmQHuksFLDF6k6ZotG9H0aILAOoCVA
rpfQuZHT6OPjoVoSMGYiRQmM+y9H9AXmvs0OwyZAoW4tNMIUV28MeBVar3TJvLwRG9uV7uVzOEhd
nAK6uqA+cf9u6K3Te6fK0tgNeGsPjssYfIbCxlBzVfk8il/E1MonRl0vtAP2p3e8l/IzoBqeOxk1
5bB4dJAwC/C6KqWGCqvWOINaoi8/MDQQOthHMEcYsjzS2kAgob1HCwXgdVQfKqpwhc7I3dvGYgBe
REp7NWejolqR3lM86ycooI6XHje9MIWFCMpbkgIZEVRejCReH39wVe37EFrj1kr7qEHCBUK5FAW7
XC3+DApwCOwrK6DU9EW7zUK04VKG3bp/Hj9yN2AI7EWDOQEYejgOcIFl5svNYdVn0fQELwWbRz2e
dAHneh45MJ/gXGY4QyxLbftRxL+/Ro63OKrp8l5ym50Uj6OJNPe6pcBJS5AtwR++VOc3JIVFPWH8
D/93CPgN//5InaTMVWYLIMBSXIwrDbNZTGCXNogTqXBNRUqDRHpvFUMKpUppJKeVPj0AIEAa2iB/
oj2NzVFELH2mRIeLIpRpZ2g6/9F2HP0rn2sL7zWeWkw7AqKEljeIC0QmZsZhUcY3FW953v0I38zQ
4+6JUsc01jaaE/F5guDDDZM8CyJdLMeaLzMksJmupXwd9DKsPhYV1is4026SjRSllgDrrPrUuuJB
UW1Meo1oDndSRik4molMqyhxWhI/WKbgHP2H5G166cxie+6lEPRR0TG0pA11+C3i+pPmmmDz0xUa
ala8YXyLIcdyIpnipPQQ9TxM10+1t3UVjtHmZLcmlyieDz/F78ZPfEdcB+TyNAJGUupIsle4A247
1TQEER3r1xBtl/1+21xEcrmBWjde6zJ7uv/JLvXTrreW7kvemJ8v2VqkXXPDPzOfeNylvBx7irK0
WR1KFKGU2yOuKbCdC58/3wn1KRe0dol3LiqxNRPQqPX6GiyOdiIoudiGdgruzIk10yiDEuXExKsQ
Qc7ma1bEqg5UrDG/zWr38v0eDcuS8y878H94dLVblHf+aOXHQOwINfS9qc2ecj5QzEd0Qz/J1mR7
YKAlsKJz7P23kltRtSPyci9KiS7tRjUuFhQd/cUq6piQN5rA+Bgda5KlOVRIEW1uia/CowuGmzsf
JxIgsZylr8f3Y5ZAWOAUTzLDguIK05lfAq3l3e4uADXV8tkR+4yFB/hAFDbtTBeDX50a1uvQ/kcV
WVX2PunCMWDBaggglb6X/iwN8Z4hO5WESfl1D4ajg/1/slYGX/ncYdcYvWpbLnRp2fgtBD2DdREo
0O4Qrm9oDQKra7RspQx3dpPGPF9j6gUCuLOOb1/LO8DNIQwu08JO1DyslauBwx++EFxJxS3WWA3F
Bl8FMO2oZJhGColDbp/aBxn19b3izbf5dMlM0UeewiwHhWzEHb0yGiTwtHbREnowa6xejXxPosD8
Uk0fw+GjQuzjqxh3PzeCiS612TGrjDejxSdIvCCCh/QtCs8KNk+x7uC6J55YN4YaIQhPSvRdUsLg
bhq2vv0UlYxSpYAeBQoyx5lcBanl8ioxjO32eN7IyVSARKgTgL1FXbEd0iUJEWA8TK1kGYBcthom
cVKFyhMU6Xa5yMTTuqnNK0E/InkOmlqYLwhWHzWNcBZtNs6YPQ4kVVNxI27gisRu33Y6Fa5beHD+
UB7sDtXP1RnvuUMr2F+XWYRGgAjIluzCJLm0WrnBawmZf/3l6hrz2qhvTiT7W2wEc+VwDAZZ3q8+
0owYxXsC7QuUBVWAXSYrZkBvisZa7tmyZGuV0beLXotNv3XbXdFdiZtKdEyMCd0dgtcNIngbtJtL
+cJ9Q18nU1BgRTJj7htGpVdD/wX0znqA0WW1vonvmNsiwdGOrDthKLwKFDDQ8S9EYvfTb8S588pc
dop8POYLrWdGE3T63aeATwf5ZY5HdfBV2cB879sV41sG2Qx/Vn52BcdFEVlXFfBZPERAbhoc9Hcq
h6NFdVoS2Zw1VsopTKqyOr6tqPh/rOrwu8Uyw3qiIQLEtdHWd6xi4k2957PuGPE/9KxKueijqNrG
/9wYsopUh/Kg3yEem0YR2vrmwYTKr9lwOpBp3F333vMhuVSUBKof5ef6hPZgvwUD14mZGu+ZxCKj
TjZNjaWFtk9E9esAiMFP5hxsIg+Dhw2DX/VupbThK5ZXNvDuN9LLC3uwfgdxY+recU6Mkl2KD42O
ln+ookzIGamP4L4rLu5UVug/9ZK5aS7z2OZSZeQJUfs3JBQoQMvuuWCVii1LoctHhBFY1FyJmfMw
UGAiFPPN6D28oEk55PitIToRpZ5TC2nPjOXl0j3D9VXaVG6jzXsANK5Z/8AQI05AeZJdDY1E9VEy
jcBH6MXkE4pZH2xmVaPCie1l8F+oJRqNHsiIK1dJkQ7X/UinY+CYYsW/BrrZUkP7xFWDQ3DQNAi6
09P2/qqeBQmij/U7mZGwhE037X+WKoEeRaPutB4uYyIQj3/ZhbPTbCqd9dmmA4MygvQhdIbocdeR
YzqWKHBdayNk0tjw9ztOcBt3eBplCvLdGovMFf+F3mV3Kqj3Uu1Z5+BfLxgXg8EZwpH+B2BN7Xex
cn4NKyR2tz4BfZYr3rtnGL4PRYSisVfAg+264Pf8tuhaRQyHgQdCg2ls9AISoqzo0WkJsFzUIIU8
uzLUWl12xE9olE4uPWqGZ5UupV9WVAHgxzX0fpbF163Oe2hWrO7qV/MtgLPO2DQxnnWXISn/KPiE
ABADLMkap9jtc8Spjg+FezyLRWRFj0huCCzI1chrflzNQDYvOcsH7fvUp4K69t8Kq/71sz5OcAHP
fpq22MX3HlzduXJW4XATGn6/YnaGo19xfWS4mFEfVOI8WBQLccGk0AA35iTXvpm2vapRD1XNJkZb
a2Fq8luqUbujy2Zxz0u10R6MvI+j1tLmIze2bISagpkevL/qJ8tQtxjlPdNjk3pqUR3sE676n3cE
1G6OFPRGrdsaU0XRI2dCM9wXtOkoMRVkf5Oi1m5KasNkDxTZIbG6ntOEmAAfir7xpiM0f9RnHUju
psO2ZfKkrUJqIjgDjmqL69TDhSQutobJhZjXU/bVjWOWbFrAK5x70HZ/sSSysxBvcroVNFOJnLRI
zYtSmm37+wcZlE4YjY97SFYSJDK1nVd0wQZPIUloYVS2In+9K8Wy9zFnN6qYaJGhxjHEp2t1jesG
IFO91olj/JJmKT0gfqkBjA9+jobXjv1jcJFDj1ij+xPTqcvf5lUGJxmDajwcaedzk7gnNdws1DXl
8+ilrbdTJL12AWhBOABbfEKm54iIf7X7i10dX/zuaDZd3AjqfDByBLOjKJMSJJD415GnxrqLtBq6
+STZGWalowRQykeYF8PpNkKIC+ca4VUpRtjdXNgBfbARgwssf7OBq15JafZOItEzTrkabpnFG9G0
tCV4b824vQ4gZo0x046bcQAi1j+thnQnmeOZlwUC+9Gl+AMIlU7efoPDzhmSNZ4a2sg3xWN/YuXc
AiU1WGS9ZuDQQfCMC+pUKBQ1uY7gsOVXyR5O0/QIKxg+8E0rv3DdJFMivu9Qu9qULo765PP0OYRG
AjyQ25y0Q8xtWWNk8iFllDxqqTNDmtTdOCklJzqU4Sp2039Wj5T4YP1dWL3Xfw7KgUrXownDau7V
yhFlfdD3oTwAdgor3PKBAjf40m6CLWABTpNj/Mt7kCdqDM2R+QLPBIWQ9UvicthxErgjf8uhiiNO
YkWHKiEykjkVzy4SJDFJF6pzckhKDwoNx2BVZE2Ed1CG8unNX4PnINtRDFIYRIKxs4BJtXhtRq3l
szYnFYO6AAwtoTlbyC9+FAk7zV7NHoRIQ6790aLQYYD0mBIU4ANqlQZg+nfN5dE71tuQkYQxBZF2
VIGNIb+n5pIrMvGnkGp4/vGj6VnTgSnXQkjOKg1GdMTCHSHMskWX9/xUQNWMYOS3GsEsxP8PnNL7
VuvR0B3u0B3bNMN5la3Bbe+pIwfWBBZsjkABlDdIfU3vqUY7/dkz/seVK+RNCQrvWoGCe4dGVVs/
xoTqeG7v6TBx5MY73cbZVz4Rwy3I7muTObtxjJQ8cjzw3aM4M8DFev5DEz8tzJDrpedkcEoOJWvh
+7awUupApIdR7waGT4Fz7WpdYTWrtJFBwWD76hE/JcMQ7J7WE/Wm2Y1Dd15aUWH3YNER42PkAhQZ
RvQoH0AuzRiUgr/m4mzoH6psNeagnGcxBnRpruSIAHY0CW47nTDJjzYe1xFPys0RTUDRej0TpVDH
W3MxztjmXYlpbkVYQdZ9KQo5DTb4CRjQWY//bJSzmQzyHf4pE4vrehC3jaLmCbZRAaH5XI3/hGZa
O7M40LNvKv2/UEJsTRPa7Z1r/W7CP3AHyVjkUm86SAG8IFt7ie6BsH5BQyLO1TQMGaRzJsH70YNE
pxY1ri0WbScsDDoZbyMugSDDglBVOAzmnqjZhJAuRPHLEL82uihYu7TXYP7O9I1rybYPphwWo0xG
Eec/REK2ryFvJeGXehozyuVozRTYLf2pLVvhSvOoyoid3GlxWRprCeT8gpSxPvcTONuAfaoKDwPn
c86h0X/S/XMJ8N5ru2gsuNBgqxdgWQ3yD3rftzOCdbtM5IAlwgZPyKtX+ohHGOVs8+lMpfrv+nJb
r6hPFJiytk6NASjB6FWJ1FUX1SAtNYz1ETUi/jYCkMu4t/H1/pb/oQlKmQOJYp9o0AxQJ0vf/ADv
/Slbvlkl0mu1sSDqW24oXS7XTWzMeqfHMRFyyevoFPwjlrrDReTdHAGNUlQpawx1wLjtLa35ZTED
nfoMM0+XKfYIVqNQuWY3ToIpu6F0vpqDwAiadnBcxdu3e5L028gt62wvPKjC0Ig5eZheshNcW/8Q
LKq/R9ekulmh244pBbDhoOqbPVdAGSRJDn8c5ifbFkqtNzG0T2RW4AmPxjVHbCo/qcPIm+8+xtuQ
qU8adJVHzq2smNeiGzq3Af+heyWzddFgv3JHAG+f1ItJ1QZNHbyzCcrB0d6GLW5DirR0rc3XuNXk
iXAKcBl//0h93V84S6my2B5XVkVNA0BW8H1QnW5KnCn4tHKlsqPaPRtPWn8xc4sFIJjeVqIRmGl8
DY5Hu7//hmd3RklN8n6KBJcFLKVx1DQpDPvjbbQs2SnPAYggRO8EdyOgDOcSr6KD/GRaqnFIwJDT
Qvvhz8q6otAljH0/P5y4unVW0IDmCiP8GtSLojOVtkuldBr8fylEr311ugA6IDfDDWkHg5jMQ29f
U2+YP7hXkc3FMKaisQnXx9nnAgV9DJ/YBGjBvHiI2cOtLzsIuSaGWdHckip3fnlSCMYEMOtgqjip
qEYh18gUC/xz/1n3PdNIwrLLecTyX5K70F25QxYogtbcTIFW6oguVwbA/ULhGAl2ODDmag1mMBoJ
VfjnNXGYyAzBuW/93GYje/HYQCFMXbm87jXl3jTJ67bDOjMTzwZLkxRHnOqkiMaCrmj4YID8Jxpn
UrNP07TiEwDkUeFyJA6agCcI9SPTyfa9MGANp5gKO5PmY+dH5iEWbFUEQMdHab/GmmWAQFnix7WX
3WjcXDWQbCTY8JuS47vtiBUby9pFVtCUXVUZYD+mWWD3K7WLeKhm8BnkpVOs93f2B4rgi6lQoLYH
UJ9KtsyMhbIiZtrNTSGOhbkilVzrCS9BeZGPiYCDVx17ua9i/ISlHZPrzLgqhLX+PFcDywkZJW4S
+bo7Ogv55kE8zg2n5nKU6jOrQjx17sUggZT7wIGkWZKTX+Gv2YhBVBhpRo/zT3VRvDt8mKe0CUJL
IVCjUDUo/Ozke12P3OvZlhaHaLkYrRi6jDo3c5c+ghBqeq+2wXcjnh0eh3ZnB5NqT1UdOwARB9+f
0M/6PZ0hN+J064jmGSgMA/HxZbOF+nRFlzWuRkWWQtrrLy6HXZa4V0tTx8sC3zUSUnQs2kr8fHmj
TGbQHTYm92MT/T7Vhs2MAE0kfoAVGePahuMHvDKqUQihU5iHOX0qqknq5HUimLFuJ8NwPPE2TNuT
Zu+1Z7X4IMJeYwWJNjA7znUKpALVgwiHUCf/NZNP72MsLNYzrA/CAeVpbfq0/LxCDPnOAJivenJp
PweGaPEB5pZdSd9XjDyqp1XVcJHiT4RazQ/xTUat8iNxATh6AO+WjEyX0hZi/kBZYj2g17s0yvws
m09lgW7XRX5+bdez6IXAYMlnFJLF1oSvzHM/ZMTVP7ti+3mWv7sFc9x2DgKQ64imCZSWFI/vnCHv
cK9yjBtt7n6S9drEhwyFe7z7+vSn4HSZSXJ5MOBQLjy+EzSpxkYnFoA41MknAhYaHwJY1s2+eD5z
dWl4U2bpCKlDtgtKr3S3uP24PZeepCIZTcqG9FNbxVfIpdMKOCSwrCjkquc/ptg6M2oVOPKVGkJj
lZrDZ+41FIHtKxmRrJLxN2+jiRUJRdMpYlYO3p9zmpg/EqRbN0gsCW6SZgpC0E2OdSFiK58DHq40
liOiMogkEDVlQsUz+PueKK95hpAKU44y/DG0XYbnQWwcqcz3x2r6E+sc8QtpjbYSrPOkSe0Q1Ivg
YvO2aWA6Qk58bFWn0pHAKdXNT11AyEd5KztDppsT+0q1Laep0vztRtubmFW1X/6/zIdoxzhaIatM
jUrwhD0kKKBr/XuMRf8Dz/kQpF9f4EzGJxgeSkQxe71/jI05Zs0KuKGxMHG6t3FgQXGvImMrJaB0
q//w+KV3QZ09O0TJUXBYwrX+pttNEtzyIGPFkWHahTUTcXMjpIc7k4GXJxnyW2MYW4UbRqpiZMuw
avesx1Z3Z6zP5PR7bPqbVE7rlaOkQsHHr+PbSp5SubLYHK+S/N0uP06Vfh5v70grvRJxvW4onoko
krVYQuG9IT73SQkI4HDN2MCK2qCFLkT+ZntzFs4UN9lo7cetYlHtxIQ7/HLCkXoPnXIph9OeMcmO
z9mQpiw9k2Ah609SD9jEGAtQ6v+y1khGrmYK7IVG0nmvuGsmtvUkbCiVgp3Gw07VADSUjyzbBV07
VgZQ3KhkvYOJaSLmyBrRWuq/lFzi1WpxvpKkEXzxVQKeqnxde9u6Q42Pnk6EoxecODKXf0Puyce7
lCAgTgTXZnojo6DzLX1osM1SpZpPUZ7V0gFfSUd7gFwo/Kd7yWG55wcIKhbSqMBPeaW4Kkt5K5fo
7kDjM6t31D8dWv+qsd12v6KWghEhPSL2bubbEQkPz58VoRS+Lt+agVUrQ/ogEdVu4vYCBFRr5Z/z
HXFMB1aJ0qF+KDfvIyDvfjVKjM1kW6H3K81TjVjNfdqfJmb+w+fnXYZp7B9KyuymLs9dnnSnDRJw
m/66RX38cNJA7SX4hH+n8e9lKZiFwk+DHwGzgnW/Qe1kzFCM7ki+Uc25kzF9pkf4dFyCHohNo6N/
LkBQsVhTN98QduFNVu8CawXpQ5RUOjdMcBm/oj9ixp1WP9+hJN74UNNMlf+covXXHPonMNaFCxOr
tgx/82jYAqR3jgwrAh+0gi4GN+dSwqkb1sBQ84rlRe55A8TtFcolJE+R1YjnF73iz6KvorctIIol
qNaJ+gQ4x2eMCSPAYXADtck69VxJU2NAZuzX1O31OvnxIGJiyW1NMgkqMsUn0mlkB8YhipFqX4Ky
JOO8StUT/attb/+DzbEKjqETxxIzSfgBZF3mfaKSaudAGE2TN7wDngmVyGeC5hGzlvU9TtwqFizz
Kbkdngia9PcSCcREr1tB6OdbzB6Eg/MaS4HV5lbKaQk891qbe71V99Zfx+/B14FjNtBUMbMdIbNe
GNJk113x70sxG0B9UMOUqIGHQ6FJuEzK+tOUYN1SNQ2PG3Rp57oRRRPJls0GrSYu3+jH4E/EYZm6
qN1as9kYqXhaqVoBEeNWw7uN7Z0xjDmqgusx4/j3XPu3XJhxrUgDldMXNfM95NyhCCRbGDdHM2sY
1a2j96fkEZYhPc+6Ww2ZZbCwS35z1E23d9jBOh1QzkPOksIl7EZ6EexACu2JS40XL7c+YGf16tVq
gEHfI1Fp5gSrWZ1JBBqhE27CO6Wqkr4QnNThgSWQ5f1I8SGWswMKY3sqaAKjUvKd7SyKovhuKyjW
DamXauYXpGf73v5+MvLNt5nudB2UTj06tOG915XDNTgL2fSmamJiezHpokfWj2/p5S6KHam6nCdQ
zXF8zjMQ/pJE5kH0tzV43LhfK3kJMcSgIVwUyUF6MpHw2sjHsoz2ZwdXXoL96M0dow1jF+zyXaue
5YG6uSAm8jFMhgqJrz6nPCVI7yj8J+GME+IoH5GBEoyTpe08OHxfkAzWmrwS4uCieoraM1uCcXxq
EXfUBUFDAWHF4fK+1w2ih3iR0QUkYoRQd4Rqz5TZMdzTiZQyfb6Y0297g8wcfxW30UEFE3OuK2eV
dLVEhLCzVIdAHPmXfq1AbHMKpJBGkiVsCciTB3F1aXeIrbUaRSeACx0GhRDxM+JG+Wm0PAohFgBK
I5tBbfyjkaJiMfabZuztAcb6J1XGIAJJbojumQbshmEtMJh3/Llt1tbTpN99T/gUEyNDp/A0t3Gi
Clbmmm5X9sHib8bsb9xWgzzWxLG4O+bCnhQmBBOhug4NSYe5uPP+KFa3ZtpcCkXU5fm2Vf7R85xm
xXgfTWhkh/VQDzfYib381pNG3F0q6qPRFhWKw+Kn7EDRjSXqAXgPV17G5bBir3zvvE8lZy4eznma
cvgDOaK8KeeAWI1Odsh9NJ7s2z9Quqg7ulGf1hSVdZahZlgdTmow/KH2OoUB7JGz2ccJEFcAQtyf
JX16uQfkhTPku0a7DfJ4BGZLrPN3SRQFnTkU4x5FJenVCve86P8RiRkjlmwX1pNSKzmJPVbXuYQ/
DJZN76UPxDepLeBoBOHtgRN90gMdVYfWlAIFRop1Hk1bMPc6ty5rxPMn/zOFIaeDP+wFq6UwIPze
OtzS7Vkqa4gDOvmTkU+aicYK6SYPQfHvPMkJIgOEV96LTp6phBEMhO8qFqEtKNEIHQaJbAqZcjd6
FxXUqJ+iQuSsPzlyh9uq0nulS3qojVWx2ul6iivFmgqbwdBJ6djwRabyq/oruw42LTuMxJe9mCBt
UqC2FC/KIzcgZ4v8au3RVmNI1MRSh+u/i5p1pSIp4gC1bSbkwpCTfAnekx0Yc/R8HK34fJB6fvFK
WsLj7DTMJYJKljSgfPXmiPB08K3qRjktO08LwFKbFT3pqENz/SMgApbgQAW5WH8sIdxKXpNzMkbF
+JE7ml3cXfdK8M+h21DVmnhKQEEBryyEPMIvRlAOj8SM7Glink8bzntBXejof7g5m2mkyVu0VtYH
f2+RreqRigFbi7TCYkJEAYL0/KCSB0XrgTZj8sm+RVgysNnSnVkLFYVxV5b8MjPKLw+Qr+SBzOG7
z1xkrewclTiR7afO8wZFm8/bHioqiL2SLh5SP0FmfZQ4mCVjG/TabccEXUbGh8w22OH5QiacXgS5
sDde4cbnonoBYNAo643NLvlg8AzmDh7Gn3a3h6b3Ze/b7Jp3y3IjAF86F6VVIuIxYy8homH73KLy
pxA9EbfxVcLfuPTSXSpXYgL8zy01sRSSLzTL1hdPZ5urtT8zxUGIbseJNI53tKYEdRdUU0R1kFMH
UGrw30Oj93Sg2tt7WEJ8bVYGuwXPG5tiGvtpE0J/U8j54CQAVm5F+6/JynZa42lTMO18ZOlVoogG
dDEOqPxSoDluLOkeGRDtyazleCZ+/tmwXKQKZqRrPqXgvDdRO7d6Iir1mQeZzzCn9VJZsIrGzXwU
ZVvqO4J0fSpxPMONbBsp+sx2cRzUUTXnpj67OtobfbrM3kMLv8zSCT4lOQi00cqzHAmz7sQw/eiQ
JlmZc5f256AhXjZO4yaCXNSqTHvmqsNfP8Y1rmj8W6nOe/8XXuFb+Dgca8BBCDkMnluhbLGf4a8o
iJJov0HJIyMV6bQa1wafIaXCm96TTSBC9D0tDMWuzLbKLKeHoI8Xg2G5UIwJZSkB1pGzOktB5BdQ
4ZGeADg1G//ytXondCQum8HwdFLgZ5dakqVmzGn6AMtK1/FEglSL25ouNX+GYcSk5X/EfQVXQPGE
vjkRvxZwDrcHC3gzFwjKHzfbyuM068BjziwH6fq1W3TBfi3psUdxys9QVBGHeQhIY/lo2UP/g9XU
Cx+WDJCcR6IpmuFGCihEByad7NW6sGbpZoELgVN9vaDvzDnTQKIxqb2W4+z3ylDkr9tIaajrhY1X
6febnR+sUtKZxfIDiNs7isoeiehJ08RLLS973MCpN0mXUvwq0KDohMNiCh3sBaNZDFdR0EJq8udA
TJXN/4EWOJnQq+5j2rNMTu9rl9SiCxNrkto7Jrnp1MthVjP3c3/WyLEFSk/ZlFM6jd2yeCsBInEI
CCAB1f/IzaygsXL5cVkw8F1B2048FO3+76ivfgp/aCEPlz0Suz4IXktaNFVmB6uCl348LTWN1Slr
s/qGhPfaJO8ZvC2BdZzMdClNbPkqHov5jv2KRTda7J+379qqDwntwRWoeEYPR04Htxlo5x9eHswP
pUCbfNXT9EruuF2Rl018tGPwxGpuV7fnwU5UWTN8rTt6wf3EIu9MhahTT5eWkpeje/Foejgr5rig
HRae0D7KC+zYhU2zMwfnE3y/SeXOAReNGbGh0h5Bh/InRUARh7R8x0J6nexwQqXMXAeswlPH6cke
gPL/QN7h2nUBnVnMT/idxxOkBdVzsl8TKlNAfH/KQbi24skG+Boe689TuowdzH4rtA6QyLLv3JGL
a5u/ko3D+ZnxIhmrJXF5ybGrnAcg5unbylLn6B+nRsh5xqZ5iJRIvL6AJIK1jMg9WqfJYkNVvGw0
QtWUfvhb/KFMZiCEMH/yaXGiNVyXL7aoVe+qt0nziPmp1IJejIbxkVZ2FzRWeDfBgeDXtM69AlqP
DJHWoSx+iWuc3Vlqiqb3/4grTQvUKx2JuuBOVoJov0Nascwq86jFpFUn4qh0hGkinkr6J85AzFYU
2VRpOe18gx6N0LSy7bPCK9F1EN3FvxQOlBaDvdaUrRJgBW+9PSBMg313Wt7+iqHW6Exu0t0lkjgK
kEVayQnqH2xxDj3uFM4DwycZYp7sc0yS5bP2hUxKnsPFlRLZGsISuYA30+57vEPBvTcXROVeu8E5
GjN1hMq4wdqicrPBchSE55xoEtvKuPZfZtZDGxfy36jf+TgNCNcavT+19dhAfGt4H4swgGhE376b
fPrOYCoZ95QZrHG0cLT7HBLnBeOfXrzbr+3ktNti7Fcxb7DoHo7Xf9vywB2eJ2Q6stUwhC/aUgRk
mB4nw6TOuOFkJCX9p54W6ETvjc6C/JXuQHEc9LNVr2nZKPzwiv2td2udnMkovnU14LRmH9pYTn2W
11TUoF6sf1/y4OTpI8MUZXYI6yDtrg+Oxs7CtA8aQEQ5O6BSPBVatHfjH/1bba0BMeE7PKwkJD/5
znJGrIy8EjOf30kWgHOHmvsO/SjTf16uhm5hweTleKYAeJYXgQf52/+CRJBT5akV5mz3w933M1IE
PHqh/0JRDv88AlZaxVyfTULqsHvZQjRTdo9Ohp9bh2PMIOYJW0L/mgwzVYEAQ1qP/dtyRMvr42O6
sBw8SKX6YGPt3Qfd8873kgpKxynMRxfY6nv3cJ4PuyYJ0Lhg6QtA0wP5pN2XKEZweUNVR+FSxwiD
i9Bz6mWiM6rwBEHKt18SE8oaa900duZ+Vaf6DZFLW8ky9nvhaL4f/lZlpReojHaMEniNhd1k4+5f
IxvyGQki8V/XPoPuEJHzcsjSAxJjXy45RMR+iDUcyPvN/8lb6fq201vyv+/ntS2aCQqWEg625cpM
Skq5dvqTG+W3wh+57ChPiKUv0RcpOC0B6T4ct/+QHnPOfx75m6Ad7zys1ij9vrg0mTulsf99jm/E
p2LgE8N/LCzphy9xuYACps3OxZ2WX+tD5wrtjudaFcZhH++Ap8VlbD7ao0LWY1P3Njr1WlsGsX+3
l4gcMEoE3FqAo5Ox/GdqL9msMqHXDWhF0sgzB4YzvQijbOyJz/v5CX3Ky5rD0/67vIwV0v7BoCgM
1Aho/BoVbCTC5uXq8tdDvWLUHkhQ4ukS0KZPRAzJF8FArnhzd0DIhbZW1ZWE8GHRAzZKuhPgN0Gb
mOapCku1x1KapJxlO8tI1nZ7mmNNEPb1QchqRp5c6r6/BPzUP+c6NVfGG5bZd7mQ3yP459SYiqeI
YQwFYz0o/O1N6np/dEwsh+BMyX2P8oZ0t5pSoEtZhGIYt1sgwbrgdRgnGkDhYUgw/MAQcDuqOOgy
tTMIO6/tkBu6TTusW52v3CAoAmgRs5KF7aGOhmT0GkT5xPmTiREZf6pP46v2Ww2zsGrYJn6VpcOF
zWlWTaqPPlgJqfX5JPaaYtDwR4DbQsJ7zDWfMWIUVJh8TKAs2VLYho6PL0+NVT7GuRNvYWUxyrPd
vX7rA290KtHM+E9Td13Z7AQJjPbtxKBXhL88Stk1ZbltAZXtxMRKAbPGTnduSezTxpFrIzwVehCJ
EPflYSVPKKXjher/c1ZRiG8DB0vc4/XZihSyVyTZm8jH+2wvp30R3FF0NC/Ysc5NWD1G24PdGMDk
Kzl5SMvm0t+wb7zTrGNnzdbZY3n4YxZ6ZbpAV8/BfOXNqM9ohX2vFv50Cy9ojcufRPKxfpCJMkRl
vF3yQJPR/M46obsY0ARxCGjl79lbXFknLxLdfDRFHYKVSVb8qmRehGE8vvCCYJaUzahaAS30PL7G
iQ8zrbcfgxYaS79nMZeEPgfJL4UVDH+Cypn+VN0JZjB3p6yqVIapLnx2a6H7LXB27nI6g3GbScMG
TveHmp12HDE7NBbcfN0n9wm2FjbdiF9hFBAGdcFTc1BbogRdAmEup1fMQ82qieIRcKNXgI2L+rxl
6d0CEtgTRwqtmcInei2OxQepqocr5BeKtDw3wumXXgdRUvqfUzTR9DO3aUiFNF/1wDpiqC7SOPHq
yCGxbDGN7jCtnVTKv9dxEysK587pZ6lIE1k+ReMAlzM0k5bR8G2fbhyvwSGSl6czoGSvYC1xW81h
VxlaAMg+eW39r8eUQhDW42udcBCnsmiGnkrXnlWsvHp9Cku60s8UR87cPH2pGiPKPqURcqZ9keoe
Z5cvqQ8d/KnDyl9NoZ3Nfrn33B8f2csjbzLKD6McUUGHzy5PSigKCu3XYebzZf/p34lVNDfenpcx
Ts+gmj+fnPEiQ3zEQmc1a+93naEfwNhbtShlNJKv/2Ovqh/zT7ompWH3u+PtsO15p32aVUWTfi8a
8aJA/aAcHcJfJYUikOmT2Eysf51N+Jyrnpf0KrEJzVAFv6fYmDcvMoe/wFq1JmVX3bIijR0/rQaQ
Vl89Znyz1LXoJI0/b7yF0Kc4CCRZThY0t0joxlFbv79Lfk9nHePckhfrpLeeEBevyPK6ayl4F2Tx
PJMYjtgjOl/EMa39XKEyBqTsiaIKlsvauK03tp2jIWi50A+zatcQ4ZuWX8arUpQMaWx/wUO2xbLs
ygZM9ySKcjqkJpmT0Rddi0VW2zlme3CdhxXKm+YNcfXQWE9h6aQvgQ1rT6lnn7QYov3kit1nY5w7
sbBCVJGaK45J7EOmggCNfMFi9tk16pWmGDuXUXTs/7kLN/ArZFWxGmXzVnBbsnkrbZPED9ZaS7sL
gv2c2J027h2ej2NoXmSRs2Ovabmq4gPt2PRKQgZojv+0TE7MQrzM7h4zTpppmpe2+I21lvuhrkfc
XeuD1uVEOD0DfAFGEEFL+PAqPcPKHsGm4RVWVlxP4XMVCpf8HjoNW/GuzFe8SwSpbwjNS4dGfkFU
OURfBCU/agjGRvsnqp0DrD1xnBuTSmLbm4oEaNNTkHEkvJKUJ23SfF2LeCj9amrCAj5uHNs3mDip
AEN4PReyfhWJIqiaOkS2zbPmdKXMSkiAvtCH9pfwvxMg6Al+I5QM+WIMkU7woCEfK6W26SSzNwFE
Guj7VY/gtAIZ1xOGUV3u/fzeeXopug7/jWsKjURVj8eS0B6fvswgJjxxoi48/QhLMRxBJ6wKZmqN
lfnyhm3XjBbeGUdF9lZ3HtGp6lnKFRavS52gciaLrDOhUXXBFC339HrSn2cAH1X6VFZqFuBQ+LIm
0d/41Dc2R2ToIfSCC1rVrWgtR/oUs6jgIRCpH+uVYb377nTlf2VfJ/W+GqtCRQhzY68cwmLZ4eLG
u0cWc9NLtlnktCsR4FYK8Aui9PjFThKIMSUxzFayz92xvHqZqIU10dBQKKpfoh1jZZUElKP4NI60
E04Vtg4NpeMhJZ3/bFaw2Mt0rvDYNCeCwE9EucYEfujgNvWKk/wI6AXmru6Wr+GpkfphlOeNvagR
yx5rT9LHQguJ3KRGNBwmsWM0UNs0IFRWjeqU6R0vS9VasqloGnBvLc6UjoNURG3XhXqc17/saMiI
b4PncldkXk+ruxscpjfVZQFo2i3RlQnAj59QYPHPbdw+qhCVUMna/erBVwCh6Fp7+YYthmMt4U4T
R1I/MPBiRwnqiknG4/WpGmmBs69mQzs+bK0R1fCjthTBdXel96p3FBkNyvOefte6LpTOz7eITCVw
nRyVc+7yMFczArclg00TbZP9E5Q2N4mtZ/4NMpXc4Z6kDKmEB2Hoi7JOyZiqDV+9aZZrFUeK7wXA
XeqjpnFjil1VNcJdbILJP9gWMKSg2cATK95RvfpF7H8ukaHavuaZPJT2dBfzXIRa7qefh+1c3rxI
iuWPaFonNJnxSAuKM8mfoAovDNGUdOLv+zUHVWHPzQvIpA5RgbbSKBSi89MWlMFGasa9VxjcII5E
F220GB9LwORmemIZv6cPc98rIFEJNcAov35wZ8rijHZv5ePAj2qOHqa7s1lm3krGpPMsYOrpHVv/
XI0ccjyfJaPpYkMpt1chS2HCb8AfEKdQNVSmb+l63J2iXZHvoDaXmNmpTRtHEsMwWkFIH+RzSWYP
qEy3ej7cpxm1ckSsSwLzCVlk5NNN2iyzWW62cZZRKWiY5Hynl9X4XZwA59OtjlXRIFSZWgqZNOPQ
TT3rYJaRzRGOnEciATj35VIAD5PBOSQoSJ587WbCNA6+nLNLjPdIdaSyAT6zKsJwhDUzvvdNgBrF
0kos1ObAjjvGr9PLC4HqUh04WIakLCRd4OIUVWNZ3cOB2+Kp0XDug8/3Jh/wuH85hX3A6hgVLNfw
fRcCunv9yP1l+rucPxLEFqV3wn5omJC4yteSQsvrTyo7K/1ac41hmIIf8Zm6NDHlaU/LrHrSHr3H
VOYPsb/bzU2shT77lL8OKSJ1g7xZ2PuMglyzkbqHEljMh2WKXT41p+6pUvcABhEG5KBaquVale3R
NzGbdV/Pgtz/t+QG4JxURj91hPr7IZoPhzXaXqjJlOPxD1KqqPEE8xojrm8ON8mzfJrzOcZRhxTW
klzegytZYr+CBCsGzWpmlzjh9Cq1ETcBoPRPPNFyw33FDVH4i8W+6LNb8n2NbZDzMjD8Q7PhgNFT
n0xZyQRWmWMH4PmuRepzMreTB2nHnivlAdsvrz4scygr1w7z7fJNuqgsxJS7PEAqw1zS3lKC4RDV
tb8vN0YM3SRoixDM8NBGv3r+04HmAE4tA/wj5QFpgvuf9XHJ4pWQhZJSYnTvdndv3MMvz4lN1/CV
q1yEzxxSM5seBpod+05nrDvsABFqtz8+wJLXJsMySUvWO9X3qtrfVoP8sFWqeUSdXqp1bsFwHr09
0XIgcgpu6MZW3uBJZxncIru4EDCw2G5UnkmkUYikHuTPLFRebJxa+WTZaeQrn/5wWZM7l7JrXftn
KiwPdo1V5tDxcUuvpnHFlJ0R+Jbg50/XW3eosjuVSQCVnwmb69FuDTKuieBhz7bv9H+Wl+SvKG2J
ya3t9YYEtHrh0Ek72m3qHSlc+73oTSigBMQiqFwphw99j73dSjMs3FzkeTKR6JCmBfWw/XwyRuKO
B7ZYekisolZD9K9B0hF1r6QVyrOF/jsylZaSFymn4wFcMftZu9nCFJx+u/LvmlwB+hYvVGMTWuY3
fSSNoH+aRi1B+m0cDK1/gklgvYwX8EDyOvG9JrZ2sWnS1KCNLKBK3ASzFz4CmSrrC/OkAIR+XNGY
XK7CGEmKDnHbJif079H+DjWbVGDXL57pWJl9JpfW4pkPjLLHfNo6x5MW9Mxiqi2GCbxUrL4B08r+
L+oSwdR9uyMUu1A61BZa20xuodAOaUtAt4rEMKnqqrqoE4+/BZtNbdzDIUsZvr97+yD5KyJJ5Vh3
RuLnK5r6S3ljSPzGbwUEGLkFs3bkmE2q5U8/DO0pEoyYVBXLhCDyYNmXCjcVaXe9wxQUHNT54pcK
3PRejUYXhqd3KnnYvdlVy/frFEAbmn3jEekwL5lKUbmB2cQaxC7yAZyyhhMqhhyLFqfLrEWq3Jg0
FQBmPSNIAUmjVtwpDR9ycJ8IFnRXk0vygtbaw6zl+/xEYMSjqg2MfC4wWsddzfbODgqHt8Ht+HgH
C3VehQl4zsGlBs7Eh+byS2PioJ5zHy3H76fl1XrO/oa5IMVJM/8ruzRlQ7MBcGTKEMLqWRBhjA28
thraQNT4B+bbAYkLQsiGrqYPlyKNr3V4fCOX6L09OAPlLpnDMHBA3qc3ABSEMHCWoNhMH9AgOKH+
4vWTyYY2hpI9o0Ba7GGDGhzZkYKyrBd2yXelJNfqRz8m6sI7jkbQlpaWaM4jZGaRkAZoEBa3Z09D
AZ8WN1Saoq+kUoihGmw/0okxfVthxPu6zIC4xrFavkJEG5OyIWk+Vbcxja7dfhi2MVT+2n1CjWtm
TQ9rcypYpwVJjXer7MWz+oUn8305lxhh0+YCWiVEztAI1Emes/5nkGFPHUmJGaoXoZ70CeZLrGbH
bDXfKS3oAzORcp5icoI/hupPZlYpWz+DZdjlsByK3OZvY8XrmCGjFsyIHa1Pzi1qdWlmFF2DXVHD
rWMStNjZbMiOlHZEFAu9BMEZ25ZEccupd6XrnVejqGnANyUcIjXyxu0o3cqAXlb3Rxe1qFOX+6lh
HR5172Xv06TvTOqPwlcgSA4JF58PnNKgSoo0gcujminj7dhJ5zaajc44esqm50LYiq72dsV8Bu88
Z+TWhPUxA0U8wI2jMIGbfRWxPKYVzKG5K9K1yFVQu1jbebJ20R764lTIu4xW/vkEBB4DUI+vHK+3
S915fKVaIcVfTjUP0/wmaV4ioQsENNNjryfnyZM+1du3sp8gU3c10WrFTlMQuTdjM+UXAXsBIaVS
/ArZpRPRb8x4IALZrp7ep/bbD3+uSv4maoSUa0g2uPizSoJidmGw1Qfmd+OQvU5KRowReQHA40kG
fnfvCcJ1O7RfzObN9Vbh7gbpJOZ/J+oIE1wZPirZiaK772/nGFzFiT4WRQGzxt2DWO60JndEu6YH
zKcZljBQ7fh+tMCVrLosGK6dHySIq8OwLOySQ+yZ+4Pp/1xn5vNLQQ24ggu+LiIY2L3JFs3cW6I2
S2dW1J9SsxyAevAcVrPC7s0Kqfzo/MveTQ7YcqFQn+BDD0Wse4qTN6d4Qd0WgeG1toQdOrdGyiTv
ZcfFwwkPE0m0HTugPRIdFb83qlAZZnYqwt5qNWDsEMvIVj+09gTjwjeCUkIafhQ0tKcFGWnfQAT1
0mfEQMKcu2gUZPydOGIAL5yfP+W1/w5qOHZPNUFZCxRBFekltBmWMwN2RVW+DVHKv9Ue0Hpda/Us
zWxSY4Qg0/7fzA1klK6hfQr7N3WIaGLZ8SDNKUXgK/mnUtkSr5ca2eaG+VCbabfpFXKGlPLNgtZW
5YWmUUIHOLq8KkK24kh8Vp3fCNgfkXL0gEMRVj0yqMRt3mjwnC2v55arugN6SuZ72w//R0U5fM+r
IiS9dHtw9U5ocP6lo1xSVy2xhmbmukoLpJx2oxLhUwd6kIFT1IfFYE8eqt9ynkC/8QRuY0yO5G1P
kTbj4u6qFwMjHbykDgRLfBmMObXcpEXr0XZNZY9I0Ec+iNP0Cod6YGfp+aMkdrNAKQlZF6vv6H2q
AF0/yTqyduwc4gzMIlVSlV/WUxMvlL4KcD/xjjsTZSB//Syia2wefyLv9dyik7OczFsdDdYbMLLz
L4ghlO+TYgwTlw8xp6+HdHt9L2+REbErROjeZmEVGOqcv4ZAGaegdm1DV8AMWNdqLnZF7CAOFHjp
gsvcrMzHeCaIiT8K0qQ99Bl3L9SlfPlG5XqGwYbYXC9b+J4QtqdQFF9G1mSS0TO0OsDH0HMKVxVZ
l82aHtGWd2c+stUWdoAQSUDG7j+xVb6r29vUMGxdnq9nIYLq9ud6Yq6ucw14YtjHQHdbFuZ787Z4
TmVnWbiiWN8VwI7lMu/tUEoW/bXwePxT4i/N8pRtrSTCCY3NcH3DQBGy7GJ+nHp3yPMIi3VBuKB+
Kob1wIXti4LbEabtRnOmQ3V82+SWyxbrOFY+ND+tlxc2iqvFXD9Tkuivo6UNt+ZDDWJqAZi+Tuv9
72gojwSsGlYTTvHNB3DX+0AnKD2s5VWnW/kTjxZmR6FrT0P9pz+sW5UpQsYCFmkTONBCrB2tGjgr
s7oxSZLrwpfhxveD0polhNo/zomzrbkd0ILKnT2bCmMY5sblrqrQV9QMXdOIifI+V5FbtruwXJbV
Yui86AuzFrobMYGMS7t2yLLUeWQQxrHD8uf8h7pMxgw36I2rfrVy37AMCNWliQzY4WgsXs1wwRW/
UV/yL3nB87ddJZWZDOqlINk9rHvxWnXfPh1co4+ceNo5CBn25ORI6q2LG9eLIrM2ACr0Ga/wXNQN
QGxxoPfX684j81A0OnV1nDlh6IQysxVzG+TMaF94jELAOYx47Y/Pe+Kv+563CY5fAxcZnVvkaDrf
iK9Z9w+7yl6rRddleWyNcFFL5pPIdcyEAqm4IGQo/c8pjyrj3xR6kaaIvpVxonZy7thWVs220rkI
bww7L6j++myk2dnjo+DIHIVMelXXo4O3lykyhB8ipVNApvTaVmMkOgFiqOZEdL5fGxGKq949JwUE
u3/Rn05yYBRh/L2z4v5gCtzR5r6ryEBP+J4eqUyKwgkDxEeP1Sj5H8vWOx3TI0GVQlJMm826vSd1
bt0QfPE+uv/eFpEKWFfYkUJfKT6lkfMu7Q2MzqiQKjH5qAiaEVDCHIZiyrqsETyo6GoiE5m6dYou
+BLa8MHKS70N+65E3z5mbrqZQzcqqTMWNis0oe/m4FP1or6UMsumsFu5+4o4l6ehiyU8PAk7lttY
ZFNKkXJmrCyoSO69it822LzHr15PrSNOPQ7egVe/suR4tWO6O+GulSRflsdUa8YfNQtmLa4fpyK9
BVuFHffsC+LQrbpCd5sXMabfyQyf3r6H1zD7FfeDoIl+WAQDPFFusNNmHDijuVlDPYhXg+t/Pc/6
HaY8tpGn1l6iXrYQoewhGTE5oRpp7ORs4Wge67QnDQcdb0EWovTXwAEAaAi1VxSYcjG4BnT1ZOkJ
c9t7iDc6Dqxm+dOanQy9NTDqz/pALsfJawDCMaHVSXYenSDhF3iJl2UhDFLVtDUe5EMRHBGANSIO
Mp2h/APBe+bHfaJNLU8AK9SvlrW2lXZ9IJeZsNTNRxPFVVga+/dwQ6LB7WVD39KvermlkksWhNEt
KGhXT+YMk0QzpzanzXuTYr0vR22tnCAhTnP6E7x4oVEzVCv0wKaKdOZKugyJ9bO6TQIv9gwd9PGD
o+N8LW6h2pNilYzVtvEJ2Wr0iRc1Ro3ROgeu+nzLl+VlOcWJIVEFwRRKZIewAw5gUaPZrjenJPAx
zVEQ/Q/qqzdvkj1Pstjlck3ooF1ORmNkjZOm0p0QAmWGiGnizoSCpJv3v7S1KQnW0zFEFN+P7f7z
bGGzfqzzoJfa/IMKkn73qt+bNbarSClcw7L5qAiYHvsuxgmpexAmjMpVVJN7SsCudjVAn3r3FfWn
saNCPuipvwYv5rkFtO0Y6VghpU75C6Bjz40kfPLK7r3vHRRuhJVwmlQbKipsbl7vNwWYM9JltBAv
h0anpIQq4ZzNNMXlEjWrDj7lRtX03Dv3YSrckYx5pPdu3D4YLSw9sBG0uSW4BEohsinOAnjvHmDE
Z+CvTO/ntztUva4LrSXKaQQrCaQo9smOUN8AQkC8PrhdzbXURkbr9kA5NggEEBEmUpVj3LhH1HY/
EVpbjaSUnmSbEw4U/ykBDTuhvNb/Wm5J95euY+ibbalFnbYiAkm1xon79Odz0XObccSoPVYqejQW
ofuXXVzZy82wUJnk3PdANZGnkToQ/1/9i5Qv/EyYLg83ehFv6lKIj9bTq6npW9Crkn2WbLPDE6B5
SUC2P9MSx5LfV/Efxy1KcauEVkUUqJpTBU9EnPHf7xTYL+zfJsDYRH7rfizrqb3tA3mkJMfupjIM
QfkhixXT476efGSVDG1aBQi8hiMXq1JzYrvnm2my2eDyNIEtVLKkknVh/14RTCBnGUTBVSQsUvjp
QfcxhwM6+cgTFqGgpJoXEBKxBQ3TeoDchudHqY6skcSsvnVQXhGzGy1Mba6Np4G6o4HOxDOmkwLd
T6JDrLSfQv/N9GJaIk9GvFJf0kDr3EdLnWFlqU1+T1Yx4s3K/QCvlJauUTQbBcLUa2swtqlPwCup
DBWS2/td0o+YCb1Jg+F8Y7u+LLduH5bG/tMKY2IhSXX9gSz1Nq/pHZBnKcaFNm6z5vdPthhoaYIf
U6OpkiHoRmoAMLdlDXm3SgAKMy5fu3208CN16vpcni1MOhJhZGdH0RPnHLiwNGB6ra68+LOrqNlo
uNrOzpx0wYU9MWXd7+Ca4okY1WRdYqyCKI5yCwqGuoTrpbSZ3XNdR9CtgaOEERYKnYtck8uBzzT0
wAHt+PMSa+tDRJDSQ7i23Edbqe3HPyElf36tYfoSCm1kIk9AVn9MduC97vU7vA68gXb9AEYzBMh7
OEn4GAw2hLgNjR4m/oOS5euEo45WmX6+fQQas8agzXwEifpZksTIprCPCGpaFGJ0YefnebgBBFbi
vCMKZ7LxzxAYNHr/UAUITH5P6KhNkrYSmjK8LfTtkyawJYVlcrsejLRKJKB7sL7QMV+b0gM4PFRa
OTNKDbCjHzcYCeJgqHGdgeY2C4HXGdys69QM4lcFAf04kKaWlC6WTbgVtjlBNsus8XgfoMRxZZSm
iod+Mhq0uYAAPuwxWHVmuq20ZJeCP6HQejixb4AVVVY3FbWuNWEBXvxl/2KsK9Nc+MAfDXI9WFAE
G8qmG+Nn4roZxhPwJftHr0MzPbHEc6ltnMX+L/xDBcbRXIqc4kXoKwROgHlT0CCHP5CV9WYXov/6
9k29biyP2hPEnp0dvXDgpFhy1yxiZX0gOfQFB+WjD1MWqRHI+kLXuUVGakuoyi5DiNsj/GcycZ3J
qe9GjpK8hJP0m91jBnwsyGp6JOp4qWoaoDt2e/3kqThBy4Ad1odxvo5wxcuDzFzIforxrTFFnkik
ioSEWDsG3Ncf+csUJ0afyuVqv5xN7FVwQwoFbL3Ul9gXcV/edV663lsyZfd8EnfVG0Cy67gTKQXP
WDpGy5lFkGEP54J1qwpsGAn3YIbMnZ2R3R+NyqEGiJSBJ4XNIz52ZaYFLixtZGFm8FvXWbUK6pOo
T4kicqrgyAiMAQhdiMWTdz3cT+6qzV1RGIvKE3vsEZ87Uoe6gdWh5YcgCWhBi5+e3LwOP5sx7bQq
XTxLZRuHNeJl2xwds6PxbtT9MsvFSe/4hTv7kOMqEyXHjwJwUbcpYR9Ri8rYSLWoZE2FmEkR9obT
bMC27+IO5lantjfUE9Qp/2wx++Cy/hjcYuWyJJY0bJBQ/K3B6NY/dyU5297p7g8+GANHKi3eOsx5
eT99ALUzuEGjZlSx3TtmaordMvym5MjTeBwM9PdLJX+Goc0HhdjEsywQocfrWSJAz45Q0t6Vhvsf
bwZM8cSzs2VbjirAAfe/nrwHq0H6mZYjz86jIaTlBNq/xnXeJcbHQoUzoQUZhZzwKFbgiHIbHcRS
zOZ8TAQUdJQmoDLsCly0asrt/Msr8W8xplcjD4Lb5ugVJPk9mEoneKlxteKYPcgfZQ04t/PHsXVL
M3mZmiODjTO3sXgP26BMsRi+cGhHFL02xSalVbm7nF47evnV/rGtWGDU3odPS6ZzDNr2vHs1HEi0
U1VG7g363Z0J1gNpT5ecNKrwrQNsEdgLvWm+Si0EVTpfeJS/T1pFDd/T35mk9vq5n1tIxUZOa07M
RQpnmThlEC+GWJVJMTyYUAcw+uEwm6maIMdBEhcRYd9rWmb2XKsXtSxjYQ1dEJS47ll7/4soqgoO
c6uEB4sL4ofZuXLwe57vf1nrKcD2Dh+0vOfFN9+F5J9c2Cz3sethYLB47YjYe0dFPRxOSvzVwIEo
//Z0KXzBVxnHCDltKSB7bSbvVjIiNB4uZlzsyXp3KrQ8Oxfa9SfGYGwKdfjKrgsEXqsIyfnZKhQz
UGTriagvghFvlLdCQ5H8nvLSqFTWULixGsThfMY6Hmq2Z3e+0p91+CWECowB7OdYyH4VYJdOdC1q
ksGeLLj5SPHhsMBDRnzAquC6hvaWv9jzm8yEp+/QHWisXW0ezwskqfzdQl7Ngq1vMJJ+nZBhUCt8
vGhvx0UoEaKCRGTJ8l4r+n7AV2Mso1TlAkVPcJemtKs6T/VvtfsUpqFCKbW9rJXWBNB03gBJRpTw
khvOs9S/x2qnWP5R3ry7XimdsUkfpZhqMkHYE95wFRYH1t3FWycu57GCEZqSPDMLExXXNd67O6Om
q33DJlaC1Y6GTAxVtCESC81KHbLF7UmYp4HzK/2zj1pYiyg2gq5TJ/DvFkCpuC6D1ITCfUPEbjbg
B7nK9LTi0Lt3VVGSFJYk5ST+SECAqjhDGEw7DXwCwRnJfalCwmh/wQ8bVeYpxL+/2P8XAheErW7R
Rs42HrcJ7g8ENst+EYOOtY2ecH1wZnCGNGDlr6tb+dVD1KGCHdO3CXZBfEXu94b1e8XyR4AP9mis
m3zLM/WRltGceLBGWKYPf2Qhfv0RdGB/NaO85VQYl7dV7MseYdTMh2KlCZe105iG6og5axcaygF6
U9tGr+z3lyErj6CdJ4VuIv09RBGpPUQU9v2DazS9UPK1C+IEs7uHCQWmikQh+dkL0LltZus02nrc
X/jCl3qGcJMbQxmWMXhRG/l3HM3Lg1Ob3ATGZvvsbHSwcNEQqsSGHb+5IbpUHyOgF9YilUzmbvvx
awm9cYTF8zLIbDBaqYuNptJnKcBXc0FooIxNLNSvAmYdmR2lcnCYrOybUiqNk7Tl5NHSJ4BhhEj+
qZKb8ktYwdoxFp1WEwCK6CP6fWf6L058eMOvc6gRi94fHCU92VKC+c3foEpKnD48RHczv3VC54Rw
WUzIONW37N+vW3W+CxYTAljg+A1Zm0DUjcL1RFOnxq4YiSiq/XQnXpUDUqJjus6sTQ/MHZvQCLce
gBnpLZ3aPHRw9UbbGmEhI/WVQJrWOA0jFhE23xhpqcV+G3DGKYc1rkomAkdRBgPYJT1uiLpZ1XQQ
f0S0ANBbixVYLfExrTp3z7LYQErJFn+9Mpz7XuX3HBUVDXGLt5RJsyg2EwaY3xB0l18sQqH0YT2P
EfJkxuqWafIKusMc0l58dP1qV4AxPqEUdUNI0+S10K0PkumMMwwgQe/mSLuD3efGgCfNhS5V9BiA
n0LrYx99Jte0DZ1/woDKwKQM8PjYuREQseKMOX83jW1AgB89MbWbxNmpLJimrADdpdCLra7rYOET
RkyeLmLtswL8ZaoE1y93rVll0bdNoZkduwz8som0H3Wzk9O/CFSGqDjzJYTsKAMb19hh6DTXdh+S
9LyU7yPJk3PIZeTkYO1cZi8B6d6yHP4J8E6slPbUcG3QE9myiGd9/y8NpRJHnbVafdEkD6XgRC4+
DGjXHCQpTvOqV6UxEFjfizcoW8UM8BuuXtWzYtUt1JwsuQzW7EmLURX42iTT1GRFAnzFyMIfh+4N
y2YFRnBe3S0P64OH09jRaRCc14mwUdnFyRXEKX2gwZTGWUkGdJDf2zZPWLKig1Cs8wR1G3kg2Y0K
j5WFP14sYYndhITfphIIRvf854+KzP7jy3qEBuIyOIUfoX+NzWl0aQUTQxL8ORl0pbVGK4ZMkCFz
ZWoTuWQlI1ZCzAPMsIoHeJfq87Au9qjTkGRU7yHLDIoQqeglkIGETVhiufwG599cgiwhgjr8LV/L
z4jFR7yFJUEBw+hOGncGSUUJ59NLhhvyTh2IIZ626I//mfqaku6NvBLLukh8kWtJHnHXkTZ+VSja
oMdOGOTPEfx+BgWEFSfoA1UufxILxRGMnPzH1GFrdwvqQWouPdxlwF6atdeXEpTTCEuj6UpaU4kJ
TSJVl6A7uBBg3TDEkQiy+hIZ6FG3RBeq41rL8ST7RhZfkDMySUJCKt/T75j/35SL8jSdmxu7+q/v
FA6AAtcr3jBxvlyCM0PgkZwwqNrYUj1SdCv4Y0M4gF6Wu3kKphthNhZV/QL7qaSczA/5lpdxLlE2
VkcNx37faDAX5kD+aOfJzoY7U62IrLjQuscu0wiZ216/9TjiQm9dy8qzEFvYvOOLoI8M0kLqXbtm
K5fF9c+5cp28rXWV7s/G3KTThlgJANsC49vmnIBwgAEgHf7Jf+bphveuopsOglpOboscsQjxRwEp
Bq6urHqJPYF3P13s27KnCPxV6lo4wHha3nWD1hh0+NZpedBqHSO6NteBuauTt4PSL1N//7SJLIIS
jw8GT01KsEy6tOFe87OASRk/vcYtc4IY9Av+QpSKsbSlYTU6D50uBHMiskBpuC/kS25nR6SBe0Ek
2R8oVqiAwt+871AODiz/WJM08mB2gScfHDtZsP7OIWSR7lAmAFFrCas/b5ewRnD3a9YXKT0+rKYc
QcrsmBua372/eUZBtscFaDfgNka3AbjyzmIaAT/oTX/Fp637HxCQS55PRrpKyH+V9YX1im5mghbZ
VKkNpqh4Be/SZOT4WP+5tXkjQz5Vy75ZgSR6I5L+yPLrru7in7pAfKbdERaRwQm+SHZWHSF99gnq
AWmd++wWlKp3Ugz4pQrl6DvceUBfYcxzi/rgH4W1oqgd5EUliVdtIRmULImojdYpyokZf2s96Jd6
uLu7EVFTxBoqJW11Xhn89QcEBQxAS/V1keJqDTxGJDAOIHIsl7FfKi00oLChn3S7AsI6kGb7RIs7
HgK/GPR1tvRoNetiEMISAo3UrNM9RlJErXAucPiaNLhsV2tEtSRV5Ryqbe6XOaI/RCoAO7d6tE5Z
+2XOIsT68wBzoQqH7XaijZ0yLRf+vCl0dfMxdsLG1uOQVFJYxwekukMS5158bUfyF3HohyZ4xZIf
+ZTRbwgaCHahMe5MoVsdcPCD8x//m93PynqC5jFgl03U2waKwu7WpjBV/0KmZxRIuEvOAicCRwc3
ZhdrCcSvWkfxZaitRM0l883JaNwkc7Y1md2Rh+O+UkytQQXztMvr2Msi/5+zn97Q7XlopljL60lo
Th+q8awxe269sdTYSRrz9GtfP+mf65IM6fyW+OFyFTyMk7rQQPYC0aIAP7v6V4WBg2D/OHuku3Yu
EUUzR4/m3ex3jsurfIRiTyySbYISHTwSIePYoSO0tjKWhrxPoBZcPHOOufbE3vM1nXuvWnprzXwo
cwMy0OWrqe4SKL9XQgA4U6UMj3oseR3lf2J3j5XKzPEyWxuq9cYKCeFlJ1xdgOCfV4rtiswP4YVj
kn7dsHPGLTZh0qHgpb6lmSCAFOKhUFtlWb07Pwxj3zbEzgTXQJNCfI7qw4/UUtEgnmJjUfl9YKYo
ar6jy60H4BgSn/9+SdiGkoc+7C+FYToQxCJseQcWyZoYNRgLkZoxHddSrhrLz8DxHxbsF4sE5SZs
noH0w5l6D5TzkNTpnRDmtMTNsu9icOBaUyOapoM/UjBoGOBwesP666jwUTGyKokcSeO3umYoXrzX
A7PM5pvzwKckEQwJumfpggxVmzDmCRxxhNof0iuhjcln2bpV1twt01mFVBS6FJg0cgYoMWH2ErWT
E2kZ9J4/fzmgPkqFIWg45Cw1xhgxb/zNsyqsmQI4ngYZnZPW7EMQRWfph8ExEP0EJsBE6KE8KcXC
sYmHLco2GlSBjVtL5NLeAzfgKlQ28hqs970=
`protect end_protected
